`timescale 1ns / 1ps

module mux1024 #(
  parameter DATA_WIDTH=16,
  parameter INDX_WIDTH=10,
  parameter ADDR_WIDTH=7
)(
  input [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] din0, din1, din2, din3, din4, din5, din6, din7, din8, din9, din10, din11, din12, din13, din14, din15, din16, din17, din18, din19, din20, din21, din22, din23, din24, din25, din26, din27, din28, din29, din30, din31, din32, din33, din34, din35, din36, din37, din38, din39, din40, din41, din42, din43, din44, din45, din46, din47, din48, din49, din50, din51, din52, din53, din54, din55, din56, din57, din58, din59, din60, din61, din62, din63, din64, din65, din66, din67, din68, din69, din70, din71, din72, din73, din74, din75, din76, din77, din78, din79, din80, din81, din82, din83, din84, din85, din86, din87, din88, din89, din90, din91, din92, din93, din94, din95, din96, din97, din98, din99, din100, din101, din102, din103, din104, din105, din106, din107, din108, din109, din110, din111, din112, din113, din114, din115, din116, din117, din118, din119, din120, din121, din122, din123, din124, din125, din126, din127, din128, din129, din130, din131, din132, din133, din134, din135, din136, din137, din138, din139, din140, din141, din142, din143, din144, din145, din146, din147, din148, din149, din150, din151, din152, din153, din154, din155, din156, din157, din158, din159, din160, din161, din162, din163, din164, din165, din166, din167, din168, din169, din170, din171, din172, din173, din174, din175, din176, din177, din178, din179, din180, din181, din182, din183, din184, din185, din186, din187, din188, din189, din190, din191, din192, din193, din194, din195, din196, din197, din198, din199, din200, din201, din202, din203, din204, din205, din206, din207, din208, din209, din210, din211, din212, din213, din214, din215, din216, din217, din218, din219, din220, din221, din222, din223, din224, din225, din226, din227, din228, din229, din230, din231, din232, din233, din234, din235, din236, din237, din238, din239, din240, din241, din242, din243, din244, din245, din246, din247, din248, din249, din250, din251, din252, din253, din254, din255, din256, din257, din258, din259, din260, din261, din262, din263, din264, din265, din266, din267, din268, din269, din270, din271, din272, din273, din274, din275, din276, din277, din278, din279, din280, din281, din282, din283, din284, din285, din286, din287, din288, din289, din290, din291, din292, din293, din294, din295, din296, din297, din298, din299, din300, din301, din302, din303, din304, din305, din306, din307, din308, din309, din310, din311, din312, din313, din314, din315, din316, din317, din318, din319, din320, din321, din322, din323, din324, din325, din326, din327, din328, din329, din330, din331, din332, din333, din334, din335, din336, din337, din338, din339, din340, din341, din342, din343, din344, din345, din346, din347, din348, din349, din350, din351, din352, din353, din354, din355, din356, din357, din358, din359, din360, din361, din362, din363, din364, din365, din366, din367, din368, din369, din370, din371, din372, din373, din374, din375, din376, din377, din378, din379, din380, din381, din382, din383, din384, din385, din386, din387, din388, din389, din390, din391, din392, din393, din394, din395, din396, din397, din398, din399, din400, din401, din402, din403, din404, din405, din406, din407, din408, din409, din410, din411, din412, din413, din414, din415, din416, din417, din418, din419, din420, din421, din422, din423, din424, din425, din426, din427, din428, din429, din430, din431, din432, din433, din434, din435, din436, din437, din438, din439, din440, din441, din442, din443, din444, din445, din446, din447, din448, din449, din450, din451, din452, din453, din454, din455, din456, din457, din458, din459, din460, din461, din462, din463, din464, din465, din466, din467, din468, din469, din470, din471, din472, din473, din474, din475, din476, din477, din478, din479, din480, din481, din482, din483, din484, din485, din486, din487, din488, din489, din490, din491, din492, din493, din494, din495, din496, din497, din498, din499, din500, din501, din502, din503, din504, din505, din506, din507, din508, din509, din510, din511, din512, din513, din514, din515, din516, din517, din518, din519, din520, din521, din522, din523, din524, din525, din526, din527, din528, din529, din530, din531, din532, din533, din534, din535, din536, din537, din538, din539, din540, din541, din542, din543, din544, din545, din546, din547, din548, din549, din550, din551, din552, din553, din554, din555, din556, din557, din558, din559, din560, din561, din562, din563, din564, din565, din566, din567, din568, din569, din570, din571, din572, din573, din574, din575, din576, din577, din578, din579, din580, din581, din582, din583, din584, din585, din586, din587, din588, din589, din590, din591, din592, din593, din594, din595, din596, din597, din598, din599, din600, din601, din602, din603, din604, din605, din606, din607, din608, din609, din610, din611, din612, din613, din614, din615, din616, din617, din618, din619, din620, din621, din622, din623, din624, din625, din626, din627, din628, din629, din630, din631, din632, din633, din634, din635, din636, din637, din638, din639, din640, din641, din642, din643, din644, din645, din646, din647, din648, din649, din650, din651, din652, din653, din654, din655, din656, din657, din658, din659, din660, din661, din662, din663, din664, din665, din666, din667, din668, din669, din670, din671, din672, din673, din674, din675, din676, din677, din678, din679, din680, din681, din682, din683, din684, din685, din686, din687, din688, din689, din690, din691, din692, din693, din694, din695, din696, din697, din698, din699, din700, din701, din702, din703, din704, din705, din706, din707, din708, din709, din710, din711, din712, din713, din714, din715, din716, din717, din718, din719, din720, din721, din722, din723, din724, din725, din726, din727, din728, din729, din730, din731, din732, din733, din734, din735, din736, din737, din738, din739, din740, din741, din742, din743, din744, din745, din746, din747, din748, din749, din750, din751, din752, din753, din754, din755, din756, din757, din758, din759, din760, din761, din762, din763, din764, din765, din766, din767, din768, din769, din770, din771, din772, din773, din774, din775, din776, din777, din778, din779, din780, din781, din782, din783, din784, din785, din786, din787, din788, din789, din790, din791, din792, din793, din794, din795, din796, din797, din798, din799, din800, din801, din802, din803, din804, din805, din806, din807, din808, din809, din810, din811, din812, din813, din814, din815, din816, din817, din818, din819, din820, din821, din822, din823, din824, din825, din826, din827, din828, din829, din830, din831, din832, din833, din834, din835, din836, din837, din838, din839, din840, din841, din842, din843, din844, din845, din846, din847, din848, din849, din850, din851, din852, din853, din854, din855, din856, din857, din858, din859, din860, din861, din862, din863, din864, din865, din866, din867, din868, din869, din870, din871, din872, din873, din874, din875, din876, din877, din878, din879, din880, din881, din882, din883, din884, din885, din886, din887, din888, din889, din890, din891, din892, din893, din894, din895, din896, din897, din898, din899, din900, din901, din902, din903, din904, din905, din906, din907, din908, din909, din910, din911, din912, din913, din914, din915, din916, din917, din918, din919, din920, din921, din922, din923, din924, din925, din926, din927, din928, din929, din930, din931, din932, din933, din934, din935, din936, din937, din938, din939, din940, din941, din942, din943, din944, din945, din946, din947, din948, din949, din950, din951, din952, din953, din954, din955, din956, din957, din958, din959, din960, din961, din962, din963, din964, din965, din966, din967, din968, din969, din970, din971, din972, din973, din974, din975, din976, din977, din978, din979, din980, din981, din982, din983, din984, din985, din986, din987, din988, din989, din990, din991, din992, din993, din994, din995, din996, din997, din998, din999, din1000, din1001, din1002, din1003, din1004, din1005, din1006, din1007, din1008, din1009, din1010, din1011, din1012, din1013, din1014, din1015, din1016, din1017, din1018, din1019, din1020, din1021, din1022, din1023,
  input [9:0] sel,
  output reg [INDX_WIDTH-1:0] indx
);

  always @(*) begin
    case(sel)
      10'd0: indx = din0[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1: indx = din1[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd2: indx = din2[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd3: indx = din3[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd4: indx = din4[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd5: indx = din5[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd6: indx = din6[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd7: indx = din7[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd8: indx = din8[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd9: indx = din9[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd10: indx = din10[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd11: indx = din11[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd12: indx = din12[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd13: indx = din13[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd14: indx = din14[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd15: indx = din15[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd16: indx = din16[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd17: indx = din17[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd18: indx = din18[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd19: indx = din19[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd20: indx = din20[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd21: indx = din21[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd22: indx = din22[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd23: indx = din23[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd24: indx = din24[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd25: indx = din25[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd26: indx = din26[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd27: indx = din27[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd28: indx = din28[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd29: indx = din29[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd30: indx = din30[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd31: indx = din31[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd32: indx = din32[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd33: indx = din33[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd34: indx = din34[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd35: indx = din35[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd36: indx = din36[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd37: indx = din37[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd38: indx = din38[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd39: indx = din39[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd40: indx = din40[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd41: indx = din41[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd42: indx = din42[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd43: indx = din43[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd44: indx = din44[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd45: indx = din45[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd46: indx = din46[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd47: indx = din47[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd48: indx = din48[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd49: indx = din49[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd50: indx = din50[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd51: indx = din51[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd52: indx = din52[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd53: indx = din53[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd54: indx = din54[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd55: indx = din55[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd56: indx = din56[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd57: indx = din57[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd58: indx = din58[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd59: indx = din59[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd60: indx = din60[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd61: indx = din61[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd62: indx = din62[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd63: indx = din63[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd64: indx = din64[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd65: indx = din65[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd66: indx = din66[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd67: indx = din67[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd68: indx = din68[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd69: indx = din69[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd70: indx = din70[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd71: indx = din71[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd72: indx = din72[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd73: indx = din73[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd74: indx = din74[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd75: indx = din75[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd76: indx = din76[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd77: indx = din77[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd78: indx = din78[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd79: indx = din79[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd80: indx = din80[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd81: indx = din81[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd82: indx = din82[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd83: indx = din83[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd84: indx = din84[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd85: indx = din85[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd86: indx = din86[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd87: indx = din87[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd88: indx = din88[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd89: indx = din89[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd90: indx = din90[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd91: indx = din91[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd92: indx = din92[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd93: indx = din93[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd94: indx = din94[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd95: indx = din95[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd96: indx = din96[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd97: indx = din97[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd98: indx = din98[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd99: indx = din99[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd100: indx = din100[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd101: indx = din101[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd102: indx = din102[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd103: indx = din103[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd104: indx = din104[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd105: indx = din105[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd106: indx = din106[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd107: indx = din107[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd108: indx = din108[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd109: indx = din109[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd110: indx = din110[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd111: indx = din111[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd112: indx = din112[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd113: indx = din113[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd114: indx = din114[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd115: indx = din115[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd116: indx = din116[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd117: indx = din117[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd118: indx = din118[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd119: indx = din119[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd120: indx = din120[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd121: indx = din121[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd122: indx = din122[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd123: indx = din123[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd124: indx = din124[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd125: indx = din125[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd126: indx = din126[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd127: indx = din127[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd128: indx = din128[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd129: indx = din129[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd130: indx = din130[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd131: indx = din131[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd132: indx = din132[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd133: indx = din133[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd134: indx = din134[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd135: indx = din135[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd136: indx = din136[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd137: indx = din137[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd138: indx = din138[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd139: indx = din139[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd140: indx = din140[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd141: indx = din141[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd142: indx = din142[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd143: indx = din143[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd144: indx = din144[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd145: indx = din145[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd146: indx = din146[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd147: indx = din147[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd148: indx = din148[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd149: indx = din149[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd150: indx = din150[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd151: indx = din151[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd152: indx = din152[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd153: indx = din153[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd154: indx = din154[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd155: indx = din155[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd156: indx = din156[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd157: indx = din157[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd158: indx = din158[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd159: indx = din159[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd160: indx = din160[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd161: indx = din161[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd162: indx = din162[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd163: indx = din163[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd164: indx = din164[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd165: indx = din165[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd166: indx = din166[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd167: indx = din167[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd168: indx = din168[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd169: indx = din169[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd170: indx = din170[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd171: indx = din171[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd172: indx = din172[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd173: indx = din173[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd174: indx = din174[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd175: indx = din175[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd176: indx = din176[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd177: indx = din177[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd178: indx = din178[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd179: indx = din179[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd180: indx = din180[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd181: indx = din181[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd182: indx = din182[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd183: indx = din183[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd184: indx = din184[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd185: indx = din185[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd186: indx = din186[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd187: indx = din187[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd188: indx = din188[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd189: indx = din189[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd190: indx = din190[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd191: indx = din191[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd192: indx = din192[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd193: indx = din193[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd194: indx = din194[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd195: indx = din195[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd196: indx = din196[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd197: indx = din197[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd198: indx = din198[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd199: indx = din199[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd200: indx = din200[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd201: indx = din201[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd202: indx = din202[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd203: indx = din203[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd204: indx = din204[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd205: indx = din205[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd206: indx = din206[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd207: indx = din207[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd208: indx = din208[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd209: indx = din209[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd210: indx = din210[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd211: indx = din211[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd212: indx = din212[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd213: indx = din213[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd214: indx = din214[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd215: indx = din215[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd216: indx = din216[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd217: indx = din217[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd218: indx = din218[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd219: indx = din219[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd220: indx = din220[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd221: indx = din221[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd222: indx = din222[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd223: indx = din223[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd224: indx = din224[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd225: indx = din225[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd226: indx = din226[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd227: indx = din227[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd228: indx = din228[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd229: indx = din229[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd230: indx = din230[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd231: indx = din231[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd232: indx = din232[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd233: indx = din233[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd234: indx = din234[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd235: indx = din235[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd236: indx = din236[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd237: indx = din237[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd238: indx = din238[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd239: indx = din239[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd240: indx = din240[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd241: indx = din241[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd242: indx = din242[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd243: indx = din243[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd244: indx = din244[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd245: indx = din245[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd246: indx = din246[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd247: indx = din247[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd248: indx = din248[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd249: indx = din249[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd250: indx = din250[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd251: indx = din251[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd252: indx = din252[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd253: indx = din253[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd254: indx = din254[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd255: indx = din255[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd256: indx = din256[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd257: indx = din257[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd258: indx = din258[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd259: indx = din259[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd260: indx = din260[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd261: indx = din261[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd262: indx = din262[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd263: indx = din263[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd264: indx = din264[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd265: indx = din265[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd266: indx = din266[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd267: indx = din267[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd268: indx = din268[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd269: indx = din269[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd270: indx = din270[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd271: indx = din271[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd272: indx = din272[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd273: indx = din273[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd274: indx = din274[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd275: indx = din275[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd276: indx = din276[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd277: indx = din277[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd278: indx = din278[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd279: indx = din279[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd280: indx = din280[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd281: indx = din281[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd282: indx = din282[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd283: indx = din283[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd284: indx = din284[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd285: indx = din285[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd286: indx = din286[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd287: indx = din287[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd288: indx = din288[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd289: indx = din289[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd290: indx = din290[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd291: indx = din291[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd292: indx = din292[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd293: indx = din293[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd294: indx = din294[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd295: indx = din295[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd296: indx = din296[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd297: indx = din297[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd298: indx = din298[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd299: indx = din299[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd300: indx = din300[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd301: indx = din301[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd302: indx = din302[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd303: indx = din303[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd304: indx = din304[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd305: indx = din305[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd306: indx = din306[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd307: indx = din307[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd308: indx = din308[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd309: indx = din309[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd310: indx = din310[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd311: indx = din311[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd312: indx = din312[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd313: indx = din313[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd314: indx = din314[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd315: indx = din315[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd316: indx = din316[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd317: indx = din317[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd318: indx = din318[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd319: indx = din319[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd320: indx = din320[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd321: indx = din321[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd322: indx = din322[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd323: indx = din323[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd324: indx = din324[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd325: indx = din325[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd326: indx = din326[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd327: indx = din327[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd328: indx = din328[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd329: indx = din329[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd330: indx = din330[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd331: indx = din331[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd332: indx = din332[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd333: indx = din333[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd334: indx = din334[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd335: indx = din335[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd336: indx = din336[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd337: indx = din337[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd338: indx = din338[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd339: indx = din339[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd340: indx = din340[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd341: indx = din341[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd342: indx = din342[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd343: indx = din343[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd344: indx = din344[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd345: indx = din345[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd346: indx = din346[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd347: indx = din347[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd348: indx = din348[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd349: indx = din349[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd350: indx = din350[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd351: indx = din351[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd352: indx = din352[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd353: indx = din353[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd354: indx = din354[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd355: indx = din355[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd356: indx = din356[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd357: indx = din357[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd358: indx = din358[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd359: indx = din359[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd360: indx = din360[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd361: indx = din361[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd362: indx = din362[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd363: indx = din363[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd364: indx = din364[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd365: indx = din365[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd366: indx = din366[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd367: indx = din367[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd368: indx = din368[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd369: indx = din369[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd370: indx = din370[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd371: indx = din371[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd372: indx = din372[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd373: indx = din373[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd374: indx = din374[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd375: indx = din375[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd376: indx = din376[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd377: indx = din377[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd378: indx = din378[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd379: indx = din379[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd380: indx = din380[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd381: indx = din381[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd382: indx = din382[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd383: indx = din383[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd384: indx = din384[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd385: indx = din385[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd386: indx = din386[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd387: indx = din387[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd388: indx = din388[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd389: indx = din389[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd390: indx = din390[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd391: indx = din391[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd392: indx = din392[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd393: indx = din393[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd394: indx = din394[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd395: indx = din395[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd396: indx = din396[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd397: indx = din397[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd398: indx = din398[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd399: indx = din399[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd400: indx = din400[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd401: indx = din401[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd402: indx = din402[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd403: indx = din403[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd404: indx = din404[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd405: indx = din405[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd406: indx = din406[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd407: indx = din407[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd408: indx = din408[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd409: indx = din409[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd410: indx = din410[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd411: indx = din411[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd412: indx = din412[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd413: indx = din413[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd414: indx = din414[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd415: indx = din415[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd416: indx = din416[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd417: indx = din417[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd418: indx = din418[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd419: indx = din419[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd420: indx = din420[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd421: indx = din421[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd422: indx = din422[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd423: indx = din423[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd424: indx = din424[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd425: indx = din425[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd426: indx = din426[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd427: indx = din427[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd428: indx = din428[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd429: indx = din429[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd430: indx = din430[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd431: indx = din431[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd432: indx = din432[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd433: indx = din433[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd434: indx = din434[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd435: indx = din435[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd436: indx = din436[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd437: indx = din437[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd438: indx = din438[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd439: indx = din439[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd440: indx = din440[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd441: indx = din441[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd442: indx = din442[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd443: indx = din443[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd444: indx = din444[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd445: indx = din445[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd446: indx = din446[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd447: indx = din447[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd448: indx = din448[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd449: indx = din449[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd450: indx = din450[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd451: indx = din451[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd452: indx = din452[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd453: indx = din453[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd454: indx = din454[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd455: indx = din455[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd456: indx = din456[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd457: indx = din457[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd458: indx = din458[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd459: indx = din459[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd460: indx = din460[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd461: indx = din461[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd462: indx = din462[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd463: indx = din463[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd464: indx = din464[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd465: indx = din465[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd466: indx = din466[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd467: indx = din467[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd468: indx = din468[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd469: indx = din469[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd470: indx = din470[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd471: indx = din471[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd472: indx = din472[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd473: indx = din473[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd474: indx = din474[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd475: indx = din475[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd476: indx = din476[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd477: indx = din477[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd478: indx = din478[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd479: indx = din479[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd480: indx = din480[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd481: indx = din481[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd482: indx = din482[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd483: indx = din483[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd484: indx = din484[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd485: indx = din485[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd486: indx = din486[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd487: indx = din487[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd488: indx = din488[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd489: indx = din489[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd490: indx = din490[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd491: indx = din491[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd492: indx = din492[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd493: indx = din493[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd494: indx = din494[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd495: indx = din495[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd496: indx = din496[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd497: indx = din497[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd498: indx = din498[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd499: indx = din499[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd500: indx = din500[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd501: indx = din501[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd502: indx = din502[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd503: indx = din503[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd504: indx = din504[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd505: indx = din505[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd506: indx = din506[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd507: indx = din507[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd508: indx = din508[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd509: indx = din509[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd510: indx = din510[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd511: indx = din511[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd512: indx = din512[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd513: indx = din513[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd514: indx = din514[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd515: indx = din515[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd516: indx = din516[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd517: indx = din517[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd518: indx = din518[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd519: indx = din519[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd520: indx = din520[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd521: indx = din521[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd522: indx = din522[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd523: indx = din523[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd524: indx = din524[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd525: indx = din525[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd526: indx = din526[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd527: indx = din527[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd528: indx = din528[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd529: indx = din529[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd530: indx = din530[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd531: indx = din531[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd532: indx = din532[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd533: indx = din533[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd534: indx = din534[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd535: indx = din535[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd536: indx = din536[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd537: indx = din537[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd538: indx = din538[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd539: indx = din539[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd540: indx = din540[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd541: indx = din541[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd542: indx = din542[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd543: indx = din543[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd544: indx = din544[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd545: indx = din545[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd546: indx = din546[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd547: indx = din547[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd548: indx = din548[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd549: indx = din549[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd550: indx = din550[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd551: indx = din551[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd552: indx = din552[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd553: indx = din553[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd554: indx = din554[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd555: indx = din555[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd556: indx = din556[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd557: indx = din557[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd558: indx = din558[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd559: indx = din559[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd560: indx = din560[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd561: indx = din561[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd562: indx = din562[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd563: indx = din563[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd564: indx = din564[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd565: indx = din565[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd566: indx = din566[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd567: indx = din567[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd568: indx = din568[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd569: indx = din569[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd570: indx = din570[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd571: indx = din571[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd572: indx = din572[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd573: indx = din573[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd574: indx = din574[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd575: indx = din575[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd576: indx = din576[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd577: indx = din577[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd578: indx = din578[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd579: indx = din579[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd580: indx = din580[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd581: indx = din581[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd582: indx = din582[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd583: indx = din583[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd584: indx = din584[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd585: indx = din585[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd586: indx = din586[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd587: indx = din587[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd588: indx = din588[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd589: indx = din589[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd590: indx = din590[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd591: indx = din591[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd592: indx = din592[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd593: indx = din593[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd594: indx = din594[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd595: indx = din595[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd596: indx = din596[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd597: indx = din597[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd598: indx = din598[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd599: indx = din599[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd600: indx = din600[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd601: indx = din601[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd602: indx = din602[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd603: indx = din603[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd604: indx = din604[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd605: indx = din605[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd606: indx = din606[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd607: indx = din607[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd608: indx = din608[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd609: indx = din609[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd610: indx = din610[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd611: indx = din611[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd612: indx = din612[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd613: indx = din613[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd614: indx = din614[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd615: indx = din615[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd616: indx = din616[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd617: indx = din617[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd618: indx = din618[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd619: indx = din619[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd620: indx = din620[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd621: indx = din621[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd622: indx = din622[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd623: indx = din623[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd624: indx = din624[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd625: indx = din625[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd626: indx = din626[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd627: indx = din627[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd628: indx = din628[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd629: indx = din629[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd630: indx = din630[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd631: indx = din631[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd632: indx = din632[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd633: indx = din633[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd634: indx = din634[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd635: indx = din635[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd636: indx = din636[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd637: indx = din637[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd638: indx = din638[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd639: indx = din639[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd640: indx = din640[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd641: indx = din641[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd642: indx = din642[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd643: indx = din643[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd644: indx = din644[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd645: indx = din645[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd646: indx = din646[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd647: indx = din647[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd648: indx = din648[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd649: indx = din649[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd650: indx = din650[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd651: indx = din651[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd652: indx = din652[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd653: indx = din653[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd654: indx = din654[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd655: indx = din655[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd656: indx = din656[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd657: indx = din657[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd658: indx = din658[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd659: indx = din659[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd660: indx = din660[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd661: indx = din661[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd662: indx = din662[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd663: indx = din663[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd664: indx = din664[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd665: indx = din665[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd666: indx = din666[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd667: indx = din667[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd668: indx = din668[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd669: indx = din669[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd670: indx = din670[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd671: indx = din671[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd672: indx = din672[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd673: indx = din673[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd674: indx = din674[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd675: indx = din675[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd676: indx = din676[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd677: indx = din677[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd678: indx = din678[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd679: indx = din679[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd680: indx = din680[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd681: indx = din681[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd682: indx = din682[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd683: indx = din683[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd684: indx = din684[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd685: indx = din685[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd686: indx = din686[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd687: indx = din687[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd688: indx = din688[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd689: indx = din689[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd690: indx = din690[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd691: indx = din691[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd692: indx = din692[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd693: indx = din693[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd694: indx = din694[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd695: indx = din695[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd696: indx = din696[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd697: indx = din697[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd698: indx = din698[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd699: indx = din699[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd700: indx = din700[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd701: indx = din701[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd702: indx = din702[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd703: indx = din703[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd704: indx = din704[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd705: indx = din705[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd706: indx = din706[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd707: indx = din707[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd708: indx = din708[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd709: indx = din709[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd710: indx = din710[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd711: indx = din711[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd712: indx = din712[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd713: indx = din713[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd714: indx = din714[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd715: indx = din715[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd716: indx = din716[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd717: indx = din717[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd718: indx = din718[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd719: indx = din719[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd720: indx = din720[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd721: indx = din721[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd722: indx = din722[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd723: indx = din723[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd724: indx = din724[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd725: indx = din725[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd726: indx = din726[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd727: indx = din727[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd728: indx = din728[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd729: indx = din729[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd730: indx = din730[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd731: indx = din731[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd732: indx = din732[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd733: indx = din733[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd734: indx = din734[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd735: indx = din735[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd736: indx = din736[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd737: indx = din737[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd738: indx = din738[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd739: indx = din739[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd740: indx = din740[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd741: indx = din741[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd742: indx = din742[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd743: indx = din743[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd744: indx = din744[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd745: indx = din745[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd746: indx = din746[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd747: indx = din747[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd748: indx = din748[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd749: indx = din749[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd750: indx = din750[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd751: indx = din751[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd752: indx = din752[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd753: indx = din753[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd754: indx = din754[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd755: indx = din755[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd756: indx = din756[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd757: indx = din757[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd758: indx = din758[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd759: indx = din759[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd760: indx = din760[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd761: indx = din761[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd762: indx = din762[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd763: indx = din763[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd764: indx = din764[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd765: indx = din765[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd766: indx = din766[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd767: indx = din767[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd768: indx = din768[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd769: indx = din769[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd770: indx = din770[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd771: indx = din771[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd772: indx = din772[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd773: indx = din773[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd774: indx = din774[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd775: indx = din775[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd776: indx = din776[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd777: indx = din777[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd778: indx = din778[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd779: indx = din779[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd780: indx = din780[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd781: indx = din781[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd782: indx = din782[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd783: indx = din783[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd784: indx = din784[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd785: indx = din785[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd786: indx = din786[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd787: indx = din787[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd788: indx = din788[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd789: indx = din789[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd790: indx = din790[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd791: indx = din791[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd792: indx = din792[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd793: indx = din793[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd794: indx = din794[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd795: indx = din795[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd796: indx = din796[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd797: indx = din797[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd798: indx = din798[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd799: indx = din799[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd800: indx = din800[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd801: indx = din801[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd802: indx = din802[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd803: indx = din803[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd804: indx = din804[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd805: indx = din805[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd806: indx = din806[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd807: indx = din807[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd808: indx = din808[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd809: indx = din809[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd810: indx = din810[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd811: indx = din811[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd812: indx = din812[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd813: indx = din813[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd814: indx = din814[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd815: indx = din815[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd816: indx = din816[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd817: indx = din817[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd818: indx = din818[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd819: indx = din819[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd820: indx = din820[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd821: indx = din821[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd822: indx = din822[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd823: indx = din823[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd824: indx = din824[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd825: indx = din825[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd826: indx = din826[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd827: indx = din827[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd828: indx = din828[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd829: indx = din829[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd830: indx = din830[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd831: indx = din831[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd832: indx = din832[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd833: indx = din833[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd834: indx = din834[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd835: indx = din835[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd836: indx = din836[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd837: indx = din837[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd838: indx = din838[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd839: indx = din839[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd840: indx = din840[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd841: indx = din841[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd842: indx = din842[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd843: indx = din843[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd844: indx = din844[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd845: indx = din845[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd846: indx = din846[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd847: indx = din847[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd848: indx = din848[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd849: indx = din849[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd850: indx = din850[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd851: indx = din851[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd852: indx = din852[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd853: indx = din853[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd854: indx = din854[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd855: indx = din855[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd856: indx = din856[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd857: indx = din857[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd858: indx = din858[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd859: indx = din859[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd860: indx = din860[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd861: indx = din861[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd862: indx = din862[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd863: indx = din863[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd864: indx = din864[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd865: indx = din865[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd866: indx = din866[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd867: indx = din867[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd868: indx = din868[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd869: indx = din869[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd870: indx = din870[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd871: indx = din871[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd872: indx = din872[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd873: indx = din873[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd874: indx = din874[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd875: indx = din875[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd876: indx = din876[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd877: indx = din877[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd878: indx = din878[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd879: indx = din879[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd880: indx = din880[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd881: indx = din881[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd882: indx = din882[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd883: indx = din883[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd884: indx = din884[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd885: indx = din885[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd886: indx = din886[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd887: indx = din887[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd888: indx = din888[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd889: indx = din889[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd890: indx = din890[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd891: indx = din891[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd892: indx = din892[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd893: indx = din893[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd894: indx = din894[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd895: indx = din895[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd896: indx = din896[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd897: indx = din897[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd898: indx = din898[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd899: indx = din899[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd900: indx = din900[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd901: indx = din901[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd902: indx = din902[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd903: indx = din903[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd904: indx = din904[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd905: indx = din905[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd906: indx = din906[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd907: indx = din907[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd908: indx = din908[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd909: indx = din909[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd910: indx = din910[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd911: indx = din911[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd912: indx = din912[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd913: indx = din913[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd914: indx = din914[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd915: indx = din915[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd916: indx = din916[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd917: indx = din917[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd918: indx = din918[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd919: indx = din919[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd920: indx = din920[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd921: indx = din921[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd922: indx = din922[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd923: indx = din923[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd924: indx = din924[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd925: indx = din925[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd926: indx = din926[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd927: indx = din927[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd928: indx = din928[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd929: indx = din929[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd930: indx = din930[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd931: indx = din931[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd932: indx = din932[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd933: indx = din933[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd934: indx = din934[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd935: indx = din935[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd936: indx = din936[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd937: indx = din937[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd938: indx = din938[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd939: indx = din939[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd940: indx = din940[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd941: indx = din941[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd942: indx = din942[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd943: indx = din943[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd944: indx = din944[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd945: indx = din945[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd946: indx = din946[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd947: indx = din947[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd948: indx = din948[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd949: indx = din949[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd950: indx = din950[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd951: indx = din951[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd952: indx = din952[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd953: indx = din953[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd954: indx = din954[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd955: indx = din955[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd956: indx = din956[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd957: indx = din957[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd958: indx = din958[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd959: indx = din959[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd960: indx = din960[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd961: indx = din961[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd962: indx = din962[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd963: indx = din963[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd964: indx = din964[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd965: indx = din965[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd966: indx = din966[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd967: indx = din967[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd968: indx = din968[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd969: indx = din969[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd970: indx = din970[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd971: indx = din971[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd972: indx = din972[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd973: indx = din973[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd974: indx = din974[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd975: indx = din975[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd976: indx = din976[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd977: indx = din977[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd978: indx = din978[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd979: indx = din979[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd980: indx = din980[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd981: indx = din981[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd982: indx = din982[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd983: indx = din983[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd984: indx = din984[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd985: indx = din985[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd986: indx = din986[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd987: indx = din987[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd988: indx = din988[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd989: indx = din989[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd990: indx = din990[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd991: indx = din991[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd992: indx = din992[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd993: indx = din993[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd994: indx = din994[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd995: indx = din995[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd996: indx = din996[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd997: indx = din997[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd998: indx = din998[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd999: indx = din999[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1000: indx = din1000[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1001: indx = din1001[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1002: indx = din1002[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1003: indx = din1003[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1004: indx = din1004[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1005: indx = din1005[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1006: indx = din1006[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1007: indx = din1007[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1008: indx = din1008[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1009: indx = din1009[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1010: indx = din1010[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1011: indx = din1011[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1012: indx = din1012[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1013: indx = din1013[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1014: indx = din1014[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1015: indx = din1015[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1016: indx = din1016[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1017: indx = din1017[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1018: indx = din1018[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1019: indx = din1019[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1020: indx = din1020[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1021: indx = din1021[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1022: indx = din1022[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      10'd1023: indx = din1023[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
    endcase
  end

endmodule

