`timescale 1ns / 1ps

module mux512 #(
  parameter DATA_WIDTH=16,
  parameter INDX_WIDTH=13,
  parameter ADDR_WIDTH=6
)(
  input [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] din0, din1, din2, din3, din4, din5, din6, din7, din8, din9, din10, din11, din12, din13, din14, din15, din16, din17, din18, din19, din20, din21, din22, din23, din24, din25, din26, din27, din28, din29, din30, din31, din32, din33, din34, din35, din36, din37, din38, din39, din40, din41, din42, din43, din44, din45, din46, din47, din48, din49, din50, din51, din52, din53, din54, din55, din56, din57, din58, din59, din60, din61, din62, din63, din64, din65, din66, din67, din68, din69, din70, din71, din72, din73, din74, din75, din76, din77, din78, din79, din80, din81, din82, din83, din84, din85, din86, din87, din88, din89, din90, din91, din92, din93, din94, din95, din96, din97, din98, din99, din100, din101, din102, din103, din104, din105, din106, din107, din108, din109, din110, din111, din112, din113, din114, din115, din116, din117, din118, din119, din120, din121, din122, din123, din124, din125, din126, din127, din128, din129, din130, din131, din132, din133, din134, din135, din136, din137, din138, din139, din140, din141, din142, din143, din144, din145, din146, din147, din148, din149, din150, din151, din152, din153, din154, din155, din156, din157, din158, din159, din160, din161, din162, din163, din164, din165, din166, din167, din168, din169, din170, din171, din172, din173, din174, din175, din176, din177, din178, din179, din180, din181, din182, din183, din184, din185, din186, din187, din188, din189, din190, din191, din192, din193, din194, din195, din196, din197, din198, din199, din200, din201, din202, din203, din204, din205, din206, din207, din208, din209, din210, din211, din212, din213, din214, din215, din216, din217, din218, din219, din220, din221, din222, din223, din224, din225, din226, din227, din228, din229, din230, din231, din232, din233, din234, din235, din236, din237, din238, din239, din240, din241, din242, din243, din244, din245, din246, din247, din248, din249, din250, din251, din252, din253, din254, din255, din256, din257, din258, din259, din260, din261, din262, din263, din264, din265, din266, din267, din268, din269, din270, din271, din272, din273, din274, din275, din276, din277, din278, din279, din280, din281, din282, din283, din284, din285, din286, din287, din288, din289, din290, din291, din292, din293, din294, din295, din296, din297, din298, din299, din300, din301, din302, din303, din304, din305, din306, din307, din308, din309, din310, din311, din312, din313, din314, din315, din316, din317, din318, din319, din320, din321, din322, din323, din324, din325, din326, din327, din328, din329, din330, din331, din332, din333, din334, din335, din336, din337, din338, din339, din340, din341, din342, din343, din344, din345, din346, din347, din348, din349, din350, din351, din352, din353, din354, din355, din356, din357, din358, din359, din360, din361, din362, din363, din364, din365, din366, din367, din368, din369, din370, din371, din372, din373, din374, din375, din376, din377, din378, din379, din380, din381, din382, din383, din384, din385, din386, din387, din388, din389, din390, din391, din392, din393, din394, din395, din396, din397, din398, din399, din400, din401, din402, din403, din404, din405, din406, din407, din408, din409, din410, din411, din412, din413, din414, din415, din416, din417, din418, din419, din420, din421, din422, din423, din424, din425, din426, din427, din428, din429, din430, din431, din432, din433, din434, din435, din436, din437, din438, din439, din440, din441, din442, din443, din444, din445, din446, din447, din448, din449, din450, din451, din452, din453, din454, din455, din456, din457, din458, din459, din460, din461, din462, din463, din464, din465, din466, din467, din468, din469, din470, din471, din472, din473, din474, din475, din476, din477, din478, din479, din480, din481, din482, din483, din484, din485, din486, din487, din488, din489, din490, din491, din492, din493, din494, din495, din496, din497, din498, din499, din500, din501, din502, din503, din504, din505, din506, din507, din508, din509, din510, din511,
  input [8:0] sel,
  output reg [INDX_WIDTH-1:0] indx
);

  always @(*) begin
    case(sel)
      9'd0: indx = din0[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd1: indx = din1[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd2: indx = din2[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd3: indx = din3[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd4: indx = din4[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd5: indx = din5[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd6: indx = din6[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd7: indx = din7[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd8: indx = din8[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd9: indx = din9[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd10: indx = din10[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd11: indx = din11[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd12: indx = din12[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd13: indx = din13[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd14: indx = din14[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd15: indx = din15[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd16: indx = din16[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd17: indx = din17[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd18: indx = din18[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd19: indx = din19[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd20: indx = din20[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd21: indx = din21[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd22: indx = din22[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd23: indx = din23[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd24: indx = din24[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd25: indx = din25[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd26: indx = din26[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd27: indx = din27[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd28: indx = din28[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd29: indx = din29[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd30: indx = din30[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd31: indx = din31[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd32: indx = din32[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd33: indx = din33[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd34: indx = din34[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd35: indx = din35[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd36: indx = din36[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd37: indx = din37[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd38: indx = din38[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd39: indx = din39[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd40: indx = din40[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd41: indx = din41[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd42: indx = din42[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd43: indx = din43[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd44: indx = din44[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd45: indx = din45[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd46: indx = din46[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd47: indx = din47[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd48: indx = din48[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd49: indx = din49[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd50: indx = din50[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd51: indx = din51[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd52: indx = din52[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd53: indx = din53[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd54: indx = din54[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd55: indx = din55[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd56: indx = din56[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd57: indx = din57[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd58: indx = din58[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd59: indx = din59[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd60: indx = din60[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd61: indx = din61[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd62: indx = din62[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd63: indx = din63[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd64: indx = din64[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd65: indx = din65[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd66: indx = din66[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd67: indx = din67[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd68: indx = din68[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd69: indx = din69[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd70: indx = din70[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd71: indx = din71[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd72: indx = din72[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd73: indx = din73[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd74: indx = din74[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd75: indx = din75[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd76: indx = din76[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd77: indx = din77[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd78: indx = din78[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd79: indx = din79[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd80: indx = din80[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd81: indx = din81[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd82: indx = din82[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd83: indx = din83[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd84: indx = din84[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd85: indx = din85[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd86: indx = din86[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd87: indx = din87[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd88: indx = din88[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd89: indx = din89[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd90: indx = din90[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd91: indx = din91[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd92: indx = din92[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd93: indx = din93[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd94: indx = din94[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd95: indx = din95[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd96: indx = din96[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd97: indx = din97[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd98: indx = din98[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd99: indx = din99[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd100: indx = din100[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd101: indx = din101[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd102: indx = din102[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd103: indx = din103[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd104: indx = din104[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd105: indx = din105[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd106: indx = din106[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd107: indx = din107[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd108: indx = din108[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd109: indx = din109[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd110: indx = din110[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd111: indx = din111[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd112: indx = din112[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd113: indx = din113[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd114: indx = din114[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd115: indx = din115[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd116: indx = din116[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd117: indx = din117[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd118: indx = din118[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd119: indx = din119[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd120: indx = din120[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd121: indx = din121[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd122: indx = din122[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd123: indx = din123[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd124: indx = din124[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd125: indx = din125[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd126: indx = din126[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd127: indx = din127[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd128: indx = din128[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd129: indx = din129[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd130: indx = din130[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd131: indx = din131[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd132: indx = din132[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd133: indx = din133[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd134: indx = din134[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd135: indx = din135[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd136: indx = din136[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd137: indx = din137[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd138: indx = din138[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd139: indx = din139[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd140: indx = din140[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd141: indx = din141[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd142: indx = din142[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd143: indx = din143[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd144: indx = din144[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd145: indx = din145[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd146: indx = din146[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd147: indx = din147[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd148: indx = din148[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd149: indx = din149[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd150: indx = din150[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd151: indx = din151[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd152: indx = din152[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd153: indx = din153[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd154: indx = din154[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd155: indx = din155[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd156: indx = din156[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd157: indx = din157[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd158: indx = din158[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd159: indx = din159[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd160: indx = din160[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd161: indx = din161[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd162: indx = din162[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd163: indx = din163[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd164: indx = din164[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd165: indx = din165[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd166: indx = din166[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd167: indx = din167[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd168: indx = din168[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd169: indx = din169[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd170: indx = din170[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd171: indx = din171[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd172: indx = din172[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd173: indx = din173[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd174: indx = din174[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd175: indx = din175[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd176: indx = din176[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd177: indx = din177[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd178: indx = din178[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd179: indx = din179[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd180: indx = din180[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd181: indx = din181[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd182: indx = din182[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd183: indx = din183[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd184: indx = din184[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd185: indx = din185[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd186: indx = din186[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd187: indx = din187[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd188: indx = din188[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd189: indx = din189[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd190: indx = din190[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd191: indx = din191[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd192: indx = din192[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd193: indx = din193[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd194: indx = din194[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd195: indx = din195[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd196: indx = din196[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd197: indx = din197[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd198: indx = din198[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd199: indx = din199[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd200: indx = din200[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd201: indx = din201[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd202: indx = din202[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd203: indx = din203[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd204: indx = din204[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd205: indx = din205[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd206: indx = din206[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd207: indx = din207[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd208: indx = din208[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd209: indx = din209[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd210: indx = din210[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd211: indx = din211[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd212: indx = din212[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd213: indx = din213[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd214: indx = din214[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd215: indx = din215[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd216: indx = din216[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd217: indx = din217[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd218: indx = din218[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd219: indx = din219[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd220: indx = din220[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd221: indx = din221[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd222: indx = din222[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd223: indx = din223[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd224: indx = din224[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd225: indx = din225[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd226: indx = din226[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd227: indx = din227[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd228: indx = din228[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd229: indx = din229[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd230: indx = din230[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd231: indx = din231[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd232: indx = din232[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd233: indx = din233[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd234: indx = din234[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd235: indx = din235[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd236: indx = din236[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd237: indx = din237[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd238: indx = din238[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd239: indx = din239[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd240: indx = din240[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd241: indx = din241[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd242: indx = din242[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd243: indx = din243[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd244: indx = din244[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd245: indx = din245[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd246: indx = din246[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd247: indx = din247[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd248: indx = din248[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd249: indx = din249[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd250: indx = din250[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd251: indx = din251[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd252: indx = din252[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd253: indx = din253[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd254: indx = din254[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd255: indx = din255[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd256: indx = din256[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd257: indx = din257[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd258: indx = din258[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd259: indx = din259[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd260: indx = din260[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd261: indx = din261[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd262: indx = din262[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd263: indx = din263[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd264: indx = din264[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd265: indx = din265[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd266: indx = din266[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd267: indx = din267[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd268: indx = din268[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd269: indx = din269[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd270: indx = din270[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd271: indx = din271[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd272: indx = din272[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd273: indx = din273[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd274: indx = din274[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd275: indx = din275[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd276: indx = din276[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd277: indx = din277[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd278: indx = din278[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd279: indx = din279[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd280: indx = din280[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd281: indx = din281[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd282: indx = din282[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd283: indx = din283[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd284: indx = din284[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd285: indx = din285[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd286: indx = din286[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd287: indx = din287[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd288: indx = din288[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd289: indx = din289[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd290: indx = din290[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd291: indx = din291[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd292: indx = din292[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd293: indx = din293[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd294: indx = din294[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd295: indx = din295[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd296: indx = din296[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd297: indx = din297[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd298: indx = din298[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd299: indx = din299[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd300: indx = din300[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd301: indx = din301[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd302: indx = din302[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd303: indx = din303[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd304: indx = din304[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd305: indx = din305[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd306: indx = din306[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd307: indx = din307[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd308: indx = din308[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd309: indx = din309[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd310: indx = din310[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd311: indx = din311[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd312: indx = din312[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd313: indx = din313[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd314: indx = din314[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd315: indx = din315[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd316: indx = din316[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd317: indx = din317[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd318: indx = din318[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd319: indx = din319[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd320: indx = din320[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd321: indx = din321[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd322: indx = din322[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd323: indx = din323[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd324: indx = din324[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd325: indx = din325[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd326: indx = din326[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd327: indx = din327[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd328: indx = din328[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd329: indx = din329[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd330: indx = din330[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd331: indx = din331[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd332: indx = din332[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd333: indx = din333[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd334: indx = din334[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd335: indx = din335[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd336: indx = din336[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd337: indx = din337[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd338: indx = din338[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd339: indx = din339[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd340: indx = din340[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd341: indx = din341[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd342: indx = din342[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd343: indx = din343[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd344: indx = din344[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd345: indx = din345[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd346: indx = din346[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd347: indx = din347[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd348: indx = din348[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd349: indx = din349[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd350: indx = din350[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd351: indx = din351[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd352: indx = din352[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd353: indx = din353[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd354: indx = din354[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd355: indx = din355[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd356: indx = din356[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd357: indx = din357[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd358: indx = din358[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd359: indx = din359[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd360: indx = din360[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd361: indx = din361[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd362: indx = din362[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd363: indx = din363[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd364: indx = din364[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd365: indx = din365[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd366: indx = din366[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd367: indx = din367[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd368: indx = din368[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd369: indx = din369[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd370: indx = din370[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd371: indx = din371[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd372: indx = din372[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd373: indx = din373[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd374: indx = din374[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd375: indx = din375[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd376: indx = din376[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd377: indx = din377[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd378: indx = din378[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd379: indx = din379[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd380: indx = din380[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd381: indx = din381[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd382: indx = din382[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd383: indx = din383[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd384: indx = din384[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd385: indx = din385[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd386: indx = din386[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd387: indx = din387[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd388: indx = din388[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd389: indx = din389[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd390: indx = din390[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd391: indx = din391[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd392: indx = din392[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd393: indx = din393[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd394: indx = din394[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd395: indx = din395[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd396: indx = din396[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd397: indx = din397[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd398: indx = din398[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd399: indx = din399[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd400: indx = din400[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd401: indx = din401[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd402: indx = din402[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd403: indx = din403[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd404: indx = din404[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd405: indx = din405[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd406: indx = din406[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd407: indx = din407[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd408: indx = din408[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd409: indx = din409[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd410: indx = din410[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd411: indx = din411[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd412: indx = din412[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd413: indx = din413[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd414: indx = din414[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd415: indx = din415[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd416: indx = din416[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd417: indx = din417[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd418: indx = din418[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd419: indx = din419[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd420: indx = din420[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd421: indx = din421[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd422: indx = din422[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd423: indx = din423[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd424: indx = din424[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd425: indx = din425[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd426: indx = din426[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd427: indx = din427[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd428: indx = din428[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd429: indx = din429[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd430: indx = din430[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd431: indx = din431[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd432: indx = din432[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd433: indx = din433[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd434: indx = din434[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd435: indx = din435[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd436: indx = din436[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd437: indx = din437[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd438: indx = din438[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd439: indx = din439[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd440: indx = din440[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd441: indx = din441[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd442: indx = din442[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd443: indx = din443[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd444: indx = din444[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd445: indx = din445[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd446: indx = din446[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd447: indx = din447[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd448: indx = din448[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd449: indx = din449[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd450: indx = din450[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd451: indx = din451[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd452: indx = din452[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd453: indx = din453[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd454: indx = din454[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd455: indx = din455[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd456: indx = din456[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd457: indx = din457[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd458: indx = din458[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd459: indx = din459[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd460: indx = din460[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd461: indx = din461[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd462: indx = din462[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd463: indx = din463[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd464: indx = din464[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd465: indx = din465[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd466: indx = din466[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd467: indx = din467[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd468: indx = din468[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd469: indx = din469[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd470: indx = din470[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd471: indx = din471[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd472: indx = din472[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd473: indx = din473[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd474: indx = din474[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd475: indx = din475[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd476: indx = din476[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd477: indx = din477[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd478: indx = din478[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd479: indx = din479[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd480: indx = din480[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd481: indx = din481[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd482: indx = din482[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd483: indx = din483[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd484: indx = din484[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd485: indx = din485[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd486: indx = din486[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd487: indx = din487[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd488: indx = din488[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd489: indx = din489[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd490: indx = din490[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd491: indx = din491[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd492: indx = din492[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd493: indx = din493[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd494: indx = din494[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd495: indx = din495[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd496: indx = din496[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd497: indx = din497[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd498: indx = din498[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd499: indx = din499[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd500: indx = din500[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd501: indx = din501[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd502: indx = din502[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd503: indx = din503[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd504: indx = din504[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd505: indx = din505[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd506: indx = din506[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd507: indx = din507[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd508: indx = din508[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd509: indx = din509[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd510: indx = din510[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
      9'd511: indx = din511[(DATA_WIDTH+INDX_WIDTH)-1:DATA_WIDTH];
    endcase
  end

endmodule

