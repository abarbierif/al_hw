`timescale 1ns / 1ps

module tb_top10();

  reg  clk;
  reg  rst_n;
  wire ready;
  reg  start;
  reg  ena;
  reg  [31:0] addra;
  reg  [255:0] dina;
  reg  [31:0] wea;
  wire [255:0] douta;
  reg  enb;
  reg  [31:0] addrb;
  reg  [31:0] dinb;
  reg  [3:0] web;
  wire [31:0] doutb;

  integer i;

  top10 dut(
    .clk(clk),
    .rst_n(rst_n),
    .ready(ready),
    .start(start),
    .clka(clk),
    .rsta(rst_n),
    .ena(ena),
    .addra(addra),
    .dina(dina),
    .wea(wea),
    .douta(douta),
    .clkb(clk),
    .rstb(rst_n),
    .enb(enb),
    .addrb(addrb),
    .dinb(dinb),
    .web(web),
    .doutb(doutb)
  );

  initial begin
    clk = 0;
    rst_n = 1;
    start = 0;

    ena = 0;
    addra = 0;
    dina = 0;
    wea = 0;

    enb = 0;
    addrb = 0;
    dinb = 0;
    web = 0;

    #10;
    rst_n=0;
    #10;
    rst_n=1;

    #10;
    ena = 1;
    wea = 32'hffffffff;
    #10

    addra = 32'd0;
    dina = {96'd0, 16'd59008, 16'd12682, 16'd9443, 16'd14055, 16'd7234, 16'd28237, 16'd47867, 16'd64693, 16'd8467, 16'd30480}; // indx = 0
    #10;
    addra = 32'd32;
    dina = {96'd0, 16'd7312, 16'd53783, 16'd48416, 16'd2954, 16'd36256, 16'd56937, 16'd42897, 16'd10385, 16'd16425, 16'd61510}; // indx = 1
    #10;
    addra = 32'd64;
    dina = {96'd0, 16'd35746, 16'd26037, 16'd50667, 16'd47390, 16'd33455, 16'd16609, 16'd33661, 16'd40649, 16'd31595, 16'd17950}; // indx = 2
    #10;
    addra = 32'd96;
    dina = {96'd0, 16'd40269, 16'd9290, 16'd1473, 16'd14133, 16'd48712, 16'd15366, 16'd57667, 16'd59049, 16'd3794, 16'd33487}; // indx = 3
    #10;
    addra = 32'd128;
    dina = {96'd0, 16'd53316, 16'd11434, 16'd11919, 16'd50555, 16'd14488, 16'd11672, 16'd17525, 16'd47199, 16'd60889, 16'd36440}; // indx = 4
    #10;
    addra = 32'd160;
    dina = {96'd0, 16'd6985, 16'd46586, 16'd1983, 16'd21036, 16'd28342, 16'd13220, 16'd1936, 16'd61743, 16'd41549, 16'd11613}; // indx = 5
    #10;
    addra = 32'd192;
    dina = {96'd0, 16'd31888, 16'd52601, 16'd45831, 16'd65435, 16'd13678, 16'd35512, 16'd40192, 16'd56596, 16'd21629, 16'd25208}; // indx = 6
    #10;
    addra = 32'd224;
    dina = {96'd0, 16'd641, 16'd56254, 16'd31699, 16'd17304, 16'd35034, 16'd26881, 16'd13630, 16'd63116, 16'd56185, 16'd18778}; // indx = 7
    #10;
    addra = 32'd256;
    dina = {96'd0, 16'd48913, 16'd18916, 16'd10221, 16'd22203, 16'd49195, 16'd60945, 16'd30903, 16'd56500, 16'd43791, 16'd14285}; // indx = 8
    #10;
    addra = 32'd288;
    dina = {96'd0, 16'd10906, 16'd28599, 16'd588, 16'd33621, 16'd48144, 16'd11091, 16'd33291, 16'd40469, 16'd53892, 16'd63781}; // indx = 9
    #10;
    addra = 32'd320;
    dina = {96'd0, 16'd64663, 16'd55951, 16'd16853, 16'd57427, 16'd20530, 16'd62494, 16'd27339, 16'd37258, 16'd9496, 16'd23625}; // indx = 10
    #10;
    addra = 32'd352;
    dina = {96'd0, 16'd39450, 16'd56026, 16'd65084, 16'd58281, 16'd29553, 16'd25015, 16'd32068, 16'd582, 16'd4033, 16'd21773}; // indx = 11
    #10;
    addra = 32'd384;
    dina = {96'd0, 16'd58631, 16'd4655, 16'd46055, 16'd34814, 16'd4119, 16'd61786, 16'd10541, 16'd15330, 16'd22976, 16'd22129}; // indx = 12
    #10;
    addra = 32'd416;
    dina = {96'd0, 16'd65440, 16'd45903, 16'd64966, 16'd14855, 16'd28349, 16'd13553, 16'd32171, 16'd65434, 16'd36953, 16'd7022}; // indx = 13
    #10;
    addra = 32'd448;
    dina = {96'd0, 16'd18343, 16'd33479, 16'd40709, 16'd50204, 16'd59587, 16'd2625, 16'd1575, 16'd12193, 16'd33647, 16'd23261}; // indx = 14
    #10;
    addra = 32'd480;
    dina = {96'd0, 16'd31416, 16'd62698, 16'd21299, 16'd41502, 16'd20898, 16'd35475, 16'd31525, 16'd37959, 16'd23739, 16'd54942}; // indx = 15
    #10;
    addra = 32'd512;
    dina = {96'd0, 16'd25643, 16'd38083, 16'd13740, 16'd34283, 16'd21873, 16'd32445, 16'd33824, 16'd7949, 16'd15460, 16'd5378}; // indx = 16
    #10;
    addra = 32'd544;
    dina = {96'd0, 16'd41543, 16'd38044, 16'd26949, 16'd40079, 16'd61775, 16'd45716, 16'd24842, 16'd42709, 16'd53857, 16'd39028}; // indx = 17
    #10;
    addra = 32'd576;
    dina = {96'd0, 16'd62767, 16'd36535, 16'd40275, 16'd33101, 16'd55068, 16'd15000, 16'd5224, 16'd7125, 16'd43927, 16'd49269}; // indx = 18
    #10;
    addra = 32'd608;
    dina = {96'd0, 16'd44099, 16'd12041, 16'd53576, 16'd27967, 16'd25534, 16'd15516, 16'd10195, 16'd36241, 16'd843, 16'd6331}; // indx = 19
    #10;
    addra = 32'd640;
    dina = {96'd0, 16'd40792, 16'd3066, 16'd31975, 16'd48297, 16'd11427, 16'd61611, 16'd34391, 16'd50790, 16'd8365, 16'd22095}; // indx = 20
    #10;
    addra = 32'd672;
    dina = {96'd0, 16'd11943, 16'd58797, 16'd46615, 16'd18296, 16'd21299, 16'd46082, 16'd3632, 16'd10776, 16'd41040, 16'd3255}; // indx = 21
    #10;
    addra = 32'd704;
    dina = {96'd0, 16'd34854, 16'd10203, 16'd15379, 16'd49650, 16'd3004, 16'd48077, 16'd65332, 16'd8697, 16'd63909, 16'd13570}; // indx = 22
    #10;
    addra = 32'd736;
    dina = {96'd0, 16'd17272, 16'd20862, 16'd41996, 16'd24839, 16'd51021, 16'd557, 16'd63226, 16'd20680, 16'd35502, 16'd40671}; // indx = 23
    #10;
    addra = 32'd768;
    dina = {96'd0, 16'd8187, 16'd53947, 16'd44328, 16'd37089, 16'd20314, 16'd17540, 16'd61732, 16'd5384, 16'd10477, 16'd45489}; // indx = 24
    #10;
    addra = 32'd800;
    dina = {96'd0, 16'd4032, 16'd31205, 16'd34708, 16'd55113, 16'd52091, 16'd25428, 16'd868, 16'd27408, 16'd34639, 16'd39346}; // indx = 25
    #10;
    addra = 32'd832;
    dina = {96'd0, 16'd12652, 16'd32736, 16'd46507, 16'd39157, 16'd13498, 16'd54010, 16'd45095, 16'd36096, 16'd49529, 16'd21768}; // indx = 26
    #10;
    addra = 32'd864;
    dina = {96'd0, 16'd39635, 16'd22309, 16'd14048, 16'd4804, 16'd7198, 16'd25276, 16'd29463, 16'd37708, 16'd52282, 16'd40316}; // indx = 27
    #10;
    addra = 32'd896;
    dina = {96'd0, 16'd42456, 16'd19689, 16'd37901, 16'd15148, 16'd2645, 16'd63153, 16'd32019, 16'd21202, 16'd24525, 16'd49849}; // indx = 28
    #10;
    addra = 32'd928;
    dina = {96'd0, 16'd35776, 16'd44231, 16'd7826, 16'd59917, 16'd33980, 16'd23199, 16'd16795, 16'd29536, 16'd40637, 16'd13909}; // indx = 29
    #10;
    addra = 32'd960;
    dina = {96'd0, 16'd27901, 16'd28788, 16'd63476, 16'd19820, 16'd55817, 16'd30331, 16'd6564, 16'd52224, 16'd40957, 16'd36412}; // indx = 30
    #10;
    addra = 32'd992;
    dina = {96'd0, 16'd13067, 16'd44209, 16'd42015, 16'd31021, 16'd10429, 16'd38931, 16'd26771, 16'd27701, 16'd33227, 16'd25707}; // indx = 31
    #10;
    addra = 32'd1024;
    dina = {96'd0, 16'd53312, 16'd18328, 16'd41857, 16'd45990, 16'd25348, 16'd61815, 16'd1551, 16'd52332, 16'd56907, 16'd61947}; // indx = 32
    #10;
    addra = 32'd1056;
    dina = {96'd0, 16'd60911, 16'd11757, 16'd35521, 16'd29239, 16'd44041, 16'd51783, 16'd53374, 16'd39066, 16'd6244, 16'd34993}; // indx = 33
    #10;
    addra = 32'd1088;
    dina = {96'd0, 16'd1324, 16'd57827, 16'd39880, 16'd20394, 16'd60287, 16'd7951, 16'd13202, 16'd50506, 16'd17519, 16'd23777}; // indx = 34
    #10;
    addra = 32'd1120;
    dina = {96'd0, 16'd18530, 16'd42002, 16'd62354, 16'd11935, 16'd32969, 16'd29399, 16'd17150, 16'd32412, 16'd63600, 16'd9771}; // indx = 35
    #10;
    addra = 32'd1152;
    dina = {96'd0, 16'd49411, 16'd21451, 16'd17525, 16'd26160, 16'd42319, 16'd33408, 16'd1619, 16'd28068, 16'd22161, 16'd53465}; // indx = 36
    #10;
    addra = 32'd1184;
    dina = {96'd0, 16'd61476, 16'd18497, 16'd33220, 16'd25713, 16'd42891, 16'd49939, 16'd3628, 16'd56819, 16'd37378, 16'd29884}; // indx = 37
    #10;
    addra = 32'd1216;
    dina = {96'd0, 16'd818, 16'd55427, 16'd54106, 16'd62875, 16'd32543, 16'd19456, 16'd28207, 16'd56662, 16'd21612, 16'd27035}; // indx = 38
    #10;
    addra = 32'd1248;
    dina = {96'd0, 16'd50308, 16'd5006, 16'd9281, 16'd65465, 16'd49833, 16'd47308, 16'd31931, 16'd18946, 16'd32097, 16'd62640}; // indx = 39
    #10;
    addra = 32'd1280;
    dina = {96'd0, 16'd61644, 16'd57454, 16'd35544, 16'd52939, 16'd58151, 16'd30268, 16'd13165, 16'd38716, 16'd11066, 16'd37754}; // indx = 40
    #10;
    addra = 32'd1312;
    dina = {96'd0, 16'd34633, 16'd17562, 16'd11394, 16'd47654, 16'd50200, 16'd3009, 16'd5939, 16'd7789, 16'd19938, 16'd16558}; // indx = 41
    #10;
    addra = 32'd1344;
    dina = {96'd0, 16'd51264, 16'd3402, 16'd9807, 16'd4466, 16'd45642, 16'd49859, 16'd6678, 16'd63516, 16'd17738, 16'd31058}; // indx = 42
    #10;
    addra = 32'd1376;
    dina = {96'd0, 16'd20713, 16'd64414, 16'd15765, 16'd57638, 16'd17974, 16'd58047, 16'd61039, 16'd26416, 16'd23847, 16'd15864}; // indx = 43
    #10;
    addra = 32'd1408;
    dina = {96'd0, 16'd8657, 16'd330, 16'd25410, 16'd19507, 16'd24474, 16'd586, 16'd37779, 16'd15518, 16'd24154, 16'd14042}; // indx = 44
    #10;
    addra = 32'd1440;
    dina = {96'd0, 16'd58734, 16'd22473, 16'd51735, 16'd40471, 16'd23646, 16'd13362, 16'd63905, 16'd17459, 16'd17039, 16'd10170}; // indx = 45
    #10;
    addra = 32'd1472;
    dina = {96'd0, 16'd33512, 16'd20869, 16'd29382, 16'd9467, 16'd25401, 16'd59141, 16'd53364, 16'd35950, 16'd28619, 16'd49158}; // indx = 46
    #10;
    addra = 32'd1504;
    dina = {96'd0, 16'd36566, 16'd45698, 16'd63994, 16'd10695, 16'd30069, 16'd58558, 16'd3765, 16'd34946, 16'd65386, 16'd53643}; // indx = 47
    #10;
    addra = 32'd1536;
    dina = {96'd0, 16'd13208, 16'd54100, 16'd43748, 16'd25754, 16'd11916, 16'd36461, 16'd25315, 16'd1049, 16'd17288, 16'd31069}; // indx = 48
    #10;
    addra = 32'd1568;
    dina = {96'd0, 16'd55591, 16'd3423, 16'd60373, 16'd28690, 16'd11361, 16'd3097, 16'd53245, 16'd44414, 16'd22527, 16'd41113}; // indx = 49
    #10;
    addra = 32'd1600;
    dina = {96'd0, 16'd42060, 16'd59873, 16'd8488, 16'd62888, 16'd37497, 16'd58474, 16'd21873, 16'd10333, 16'd18497, 16'd51798}; // indx = 50
    #10;
    addra = 32'd1632;
    dina = {96'd0, 16'd9767, 16'd28644, 16'd63544, 16'd46024, 16'd61010, 16'd2240, 16'd9689, 16'd20618, 16'd161, 16'd4743}; // indx = 51
    #10;
    addra = 32'd1664;
    dina = {96'd0, 16'd37037, 16'd38069, 16'd10722, 16'd63514, 16'd49557, 16'd55573, 16'd17291, 16'd46251, 16'd5968, 16'd37969}; // indx = 52
    #10;
    addra = 32'd1696;
    dina = {96'd0, 16'd26324, 16'd22388, 16'd7868, 16'd19311, 16'd25979, 16'd38277, 16'd65491, 16'd25183, 16'd9215, 16'd46474}; // indx = 53
    #10;
    addra = 32'd1728;
    dina = {96'd0, 16'd19377, 16'd49716, 16'd37692, 16'd57375, 16'd56004, 16'd32027, 16'd60840, 16'd1177, 16'd10348, 16'd58367}; // indx = 54
    #10;
    addra = 32'd1760;
    dina = {96'd0, 16'd15076, 16'd31269, 16'd22314, 16'd23680, 16'd48790, 16'd53766, 16'd43871, 16'd24418, 16'd24130, 16'd23800}; // indx = 55
    #10;
    addra = 32'd1792;
    dina = {96'd0, 16'd4529, 16'd30648, 16'd8909, 16'd60809, 16'd12945, 16'd58058, 16'd60364, 16'd19015, 16'd29949, 16'd1040}; // indx = 56
    #10;
    addra = 32'd1824;
    dina = {96'd0, 16'd6423, 16'd54464, 16'd13288, 16'd31549, 16'd38482, 16'd2831, 16'd2038, 16'd44522, 16'd57322, 16'd45013}; // indx = 57
    #10;
    addra = 32'd1856;
    dina = {96'd0, 16'd25768, 16'd63421, 16'd45379, 16'd29012, 16'd25659, 16'd63839, 16'd21501, 16'd42437, 16'd9707, 16'd63477}; // indx = 58
    #10;
    addra = 32'd1888;
    dina = {96'd0, 16'd19000, 16'd24398, 16'd28145, 16'd46040, 16'd44381, 16'd12871, 16'd64521, 16'd43261, 16'd33130, 16'd54010}; // indx = 59
    #10;
    addra = 32'd1920;
    dina = {96'd0, 16'd63037, 16'd45109, 16'd55360, 16'd8438, 16'd28303, 16'd6176, 16'd53177, 16'd63138, 16'd65172, 16'd19698}; // indx = 60
    #10;
    addra = 32'd1952;
    dina = {96'd0, 16'd34540, 16'd58185, 16'd28732, 16'd1134, 16'd21779, 16'd13618, 16'd63271, 16'd24143, 16'd61121, 16'd53957}; // indx = 61
    #10;
    addra = 32'd1984;
    dina = {96'd0, 16'd17275, 16'd14376, 16'd3964, 16'd59855, 16'd15961, 16'd26210, 16'd27466, 16'd46153, 16'd12712, 16'd38440}; // indx = 62
    #10;
    addra = 32'd2016;
    dina = {96'd0, 16'd12395, 16'd19870, 16'd55327, 16'd14774, 16'd22764, 16'd17070, 16'd47909, 16'd31001, 16'd34306, 16'd1992}; // indx = 63
    #10;
    addra = 32'd2048;
    dina = {96'd0, 16'd15576, 16'd30218, 16'd65242, 16'd23860, 16'd54331, 16'd21676, 16'd9697, 16'd34706, 16'd36980, 16'd31730}; // indx = 64
    #10;
    addra = 32'd2080;
    dina = {96'd0, 16'd6041, 16'd59484, 16'd54119, 16'd19944, 16'd9457, 16'd29214, 16'd60098, 16'd62086, 16'd21644, 16'd4482}; // indx = 65
    #10;
    addra = 32'd2112;
    dina = {96'd0, 16'd63076, 16'd26950, 16'd46610, 16'd31165, 16'd48923, 16'd29733, 16'd17046, 16'd41245, 16'd38844, 16'd39869}; // indx = 66
    #10;
    addra = 32'd2144;
    dina = {96'd0, 16'd54424, 16'd47279, 16'd24755, 16'd51386, 16'd30577, 16'd61933, 16'd23734, 16'd39586, 16'd35228, 16'd30922}; // indx = 67
    #10;
    addra = 32'd2176;
    dina = {96'd0, 16'd54042, 16'd44831, 16'd53466, 16'd52006, 16'd56103, 16'd24549, 16'd7565, 16'd4272, 16'd25173, 16'd34630}; // indx = 68
    #10;
    addra = 32'd2208;
    dina = {96'd0, 16'd24341, 16'd25827, 16'd59281, 16'd58374, 16'd54363, 16'd58747, 16'd18767, 16'd42901, 16'd18579, 16'd16419}; // indx = 69
    #10;
    addra = 32'd2240;
    dina = {96'd0, 16'd47926, 16'd16167, 16'd16331, 16'd2122, 16'd54186, 16'd40083, 16'd21001, 16'd3941, 16'd7056, 16'd29431}; // indx = 70
    #10;
    addra = 32'd2272;
    dina = {96'd0, 16'd41803, 16'd65267, 16'd60656, 16'd2511, 16'd15667, 16'd39560, 16'd20705, 16'd51495, 16'd11091, 16'd25243}; // indx = 71
    #10;
    addra = 32'd2304;
    dina = {96'd0, 16'd17942, 16'd10368, 16'd3461, 16'd23226, 16'd65451, 16'd35105, 16'd51890, 16'd41534, 16'd43628, 16'd47637}; // indx = 72
    #10;
    addra = 32'd2336;
    dina = {96'd0, 16'd8167, 16'd27334, 16'd36036, 16'd49713, 16'd31708, 16'd6161, 16'd25482, 16'd15323, 16'd27672, 16'd42261}; // indx = 73
    #10;
    addra = 32'd2368;
    dina = {96'd0, 16'd53277, 16'd2605, 16'd25486, 16'd18745, 16'd44483, 16'd48342, 16'd59634, 16'd12082, 16'd6838, 16'd35646}; // indx = 74
    #10;
    addra = 32'd2400;
    dina = {96'd0, 16'd51569, 16'd31783, 16'd48021, 16'd53549, 16'd42031, 16'd35431, 16'd19852, 16'd9418, 16'd33939, 16'd26372}; // indx = 75
    #10;
    addra = 32'd2432;
    dina = {96'd0, 16'd15098, 16'd30789, 16'd3661, 16'd58231, 16'd51329, 16'd34525, 16'd10616, 16'd7760, 16'd19762, 16'd57264}; // indx = 76
    #10;
    addra = 32'd2464;
    dina = {96'd0, 16'd32152, 16'd61880, 16'd57007, 16'd61647, 16'd8118, 16'd50395, 16'd18461, 16'd7819, 16'd16246, 16'd55465}; // indx = 77
    #10;
    addra = 32'd2496;
    dina = {96'd0, 16'd58758, 16'd25804, 16'd8798, 16'd39428, 16'd4789, 16'd24282, 16'd55063, 16'd43848, 16'd17803, 16'd2081}; // indx = 78
    #10;
    addra = 32'd2528;
    dina = {96'd0, 16'd57424, 16'd57680, 16'd7763, 16'd65366, 16'd2955, 16'd305, 16'd29697, 16'd17466, 16'd48280, 16'd2600}; // indx = 79
    #10;
    addra = 32'd2560;
    dina = {96'd0, 16'd7141, 16'd45852, 16'd54982, 16'd45003, 16'd39479, 16'd64397, 16'd31401, 16'd45053, 16'd43858, 16'd53470}; // indx = 80
    #10;
    addra = 32'd2592;
    dina = {96'd0, 16'd27132, 16'd5651, 16'd63481, 16'd57430, 16'd14942, 16'd64909, 16'd41964, 16'd53293, 16'd31188, 16'd11860}; // indx = 81
    #10;
    addra = 32'd2624;
    dina = {96'd0, 16'd21274, 16'd6563, 16'd28346, 16'd52633, 16'd56364, 16'd28550, 16'd48183, 16'd35647, 16'd16104, 16'd39981}; // indx = 82
    #10;
    addra = 32'd2656;
    dina = {96'd0, 16'd23937, 16'd59983, 16'd17202, 16'd31531, 16'd62404, 16'd27474, 16'd53075, 16'd22883, 16'd14768, 16'd25496}; // indx = 83
    #10;
    addra = 32'd2688;
    dina = {96'd0, 16'd10768, 16'd3273, 16'd11602, 16'd57226, 16'd2981, 16'd2047, 16'd55609, 16'd24837, 16'd42829, 16'd52320}; // indx = 84
    #10;
    addra = 32'd2720;
    dina = {96'd0, 16'd50904, 16'd59941, 16'd10195, 16'd42460, 16'd56406, 16'd39843, 16'd24658, 16'd21419, 16'd32825, 16'd21401}; // indx = 85
    #10;
    addra = 32'd2752;
    dina = {96'd0, 16'd51125, 16'd47325, 16'd46966, 16'd18683, 16'd28996, 16'd61634, 16'd62026, 16'd64767, 16'd50106, 16'd22114}; // indx = 86
    #10;
    addra = 32'd2784;
    dina = {96'd0, 16'd7022, 16'd28236, 16'd25987, 16'd50161, 16'd41426, 16'd52555, 16'd17524, 16'd40546, 16'd18355, 16'd53793}; // indx = 87
    #10;
    addra = 32'd2816;
    dina = {96'd0, 16'd14893, 16'd62378, 16'd54396, 16'd19356, 16'd50443, 16'd50576, 16'd37111, 16'd54352, 16'd33565, 16'd31701}; // indx = 88
    #10;
    addra = 32'd2848;
    dina = {96'd0, 16'd54046, 16'd32066, 16'd58706, 16'd13841, 16'd12677, 16'd8544, 16'd45709, 16'd60123, 16'd55967, 16'd65141}; // indx = 89
    #10;
    addra = 32'd2880;
    dina = {96'd0, 16'd3281, 16'd47450, 16'd7320, 16'd57764, 16'd20028, 16'd54693, 16'd50030, 16'd26193, 16'd30772, 16'd47730}; // indx = 90
    #10;
    addra = 32'd2912;
    dina = {96'd0, 16'd22923, 16'd28965, 16'd2248, 16'd55339, 16'd59452, 16'd6029, 16'd51555, 16'd28590, 16'd32728, 16'd57514}; // indx = 91
    #10;
    addra = 32'd2944;
    dina = {96'd0, 16'd9673, 16'd53890, 16'd51303, 16'd9874, 16'd54054, 16'd48088, 16'd25638, 16'd24284, 16'd61404, 16'd16061}; // indx = 92
    #10;
    addra = 32'd2976;
    dina = {96'd0, 16'd22442, 16'd13107, 16'd18450, 16'd45954, 16'd6227, 16'd4184, 16'd49509, 16'd50216, 16'd29597, 16'd29329}; // indx = 93
    #10;
    addra = 32'd3008;
    dina = {96'd0, 16'd5942, 16'd51811, 16'd40069, 16'd56710, 16'd30831, 16'd51904, 16'd30950, 16'd16183, 16'd36823, 16'd40301}; // indx = 94
    #10;
    addra = 32'd3040;
    dina = {96'd0, 16'd3348, 16'd23880, 16'd59003, 16'd12649, 16'd63817, 16'd23126, 16'd19963, 16'd5448, 16'd57836, 16'd55814}; // indx = 95
    #10;
    addra = 32'd3072;
    dina = {96'd0, 16'd57835, 16'd63908, 16'd29638, 16'd42484, 16'd45517, 16'd51688, 16'd1446, 16'd53950, 16'd55369, 16'd37518}; // indx = 96
    #10;
    addra = 32'd3104;
    dina = {96'd0, 16'd55895, 16'd34877, 16'd13392, 16'd16374, 16'd37568, 16'd48494, 16'd63204, 16'd3022, 16'd9302, 16'd17628}; // indx = 97
    #10;
    addra = 32'd3136;
    dina = {96'd0, 16'd5087, 16'd40708, 16'd46941, 16'd31187, 16'd5527, 16'd33715, 16'd11287, 16'd56497, 16'd24594, 16'd31130}; // indx = 98
    #10;
    addra = 32'd3168;
    dina = {96'd0, 16'd48165, 16'd49903, 16'd596, 16'd42245, 16'd21046, 16'd64600, 16'd13171, 16'd43497, 16'd48601, 16'd18774}; // indx = 99
    #10;
    addra = 32'd3200;
    dina = {96'd0, 16'd22115, 16'd20006, 16'd44346, 16'd53201, 16'd49682, 16'd45385, 16'd22270, 16'd39697, 16'd31954, 16'd64228}; // indx = 100
    #10;
    addra = 32'd3232;
    dina = {96'd0, 16'd32083, 16'd30957, 16'd33213, 16'd141, 16'd34469, 16'd18669, 16'd26407, 16'd41586, 16'd3255, 16'd19098}; // indx = 101
    #10;
    addra = 32'd3264;
    dina = {96'd0, 16'd6862, 16'd52274, 16'd33388, 16'd48195, 16'd43096, 16'd55831, 16'd27577, 16'd61780, 16'd19261, 16'd6835}; // indx = 102
    #10;
    addra = 32'd3296;
    dina = {96'd0, 16'd50831, 16'd42577, 16'd54561, 16'd22658, 16'd55044, 16'd11930, 16'd60972, 16'd61698, 16'd28132, 16'd41853}; // indx = 103
    #10;
    addra = 32'd3328;
    dina = {96'd0, 16'd55572, 16'd55543, 16'd27148, 16'd738, 16'd60806, 16'd33334, 16'd33257, 16'd31206, 16'd10193, 16'd16497}; // indx = 104
    #10;
    addra = 32'd3360;
    dina = {96'd0, 16'd64618, 16'd46348, 16'd35116, 16'd33470, 16'd9589, 16'd3596, 16'd30794, 16'd49128, 16'd56133, 16'd47091}; // indx = 105
    #10;
    addra = 32'd3392;
    dina = {96'd0, 16'd28894, 16'd23783, 16'd64859, 16'd43638, 16'd57008, 16'd325, 16'd51616, 16'd19427, 16'd3043, 16'd60125}; // indx = 106
    #10;
    addra = 32'd3424;
    dina = {96'd0, 16'd49639, 16'd6197, 16'd17513, 16'd37893, 16'd48719, 16'd46617, 16'd60668, 16'd116, 16'd22948, 16'd33016}; // indx = 107
    #10;
    addra = 32'd3456;
    dina = {96'd0, 16'd28311, 16'd3842, 16'd62432, 16'd12860, 16'd55081, 16'd40809, 16'd34471, 16'd4108, 16'd35957, 16'd22878}; // indx = 108
    #10;
    addra = 32'd3488;
    dina = {96'd0, 16'd42332, 16'd11327, 16'd9239, 16'd6656, 16'd55446, 16'd5055, 16'd55906, 16'd31649, 16'd24731, 16'd56297}; // indx = 109
    #10;
    addra = 32'd3520;
    dina = {96'd0, 16'd50191, 16'd53383, 16'd31905, 16'd37464, 16'd10642, 16'd31410, 16'd48313, 16'd6829, 16'd55541, 16'd24271}; // indx = 110
    #10;
    addra = 32'd3552;
    dina = {96'd0, 16'd61150, 16'd23494, 16'd59282, 16'd33764, 16'd26431, 16'd27970, 16'd52409, 16'd56395, 16'd43055, 16'd31836}; // indx = 111
    #10;
    addra = 32'd3584;
    dina = {96'd0, 16'd48394, 16'd54995, 16'd48225, 16'd10229, 16'd49209, 16'd53710, 16'd2561, 16'd35461, 16'd27574, 16'd25655}; // indx = 112
    #10;
    addra = 32'd3616;
    dina = {96'd0, 16'd41390, 16'd28104, 16'd49315, 16'd23250, 16'd52850, 16'd47659, 16'd60376, 16'd64193, 16'd22007, 16'd63976}; // indx = 113
    #10;
    addra = 32'd3648;
    dina = {96'd0, 16'd63962, 16'd10843, 16'd31804, 16'd22231, 16'd35997, 16'd10964, 16'd63971, 16'd23261, 16'd33694, 16'd59490}; // indx = 114
    #10;
    addra = 32'd3680;
    dina = {96'd0, 16'd28213, 16'd63047, 16'd52496, 16'd44927, 16'd34894, 16'd33678, 16'd16355, 16'd39908, 16'd29726, 16'd11933}; // indx = 115
    #10;
    addra = 32'd3712;
    dina = {96'd0, 16'd38341, 16'd35708, 16'd37423, 16'd25692, 16'd58905, 16'd11535, 16'd27353, 16'd58806, 16'd8646, 16'd60274}; // indx = 116
    #10;
    addra = 32'd3744;
    dina = {96'd0, 16'd44920, 16'd39591, 16'd17454, 16'd27847, 16'd15321, 16'd64629, 16'd52363, 16'd58999, 16'd49864, 16'd46112}; // indx = 117
    #10;
    addra = 32'd3776;
    dina = {96'd0, 16'd50299, 16'd39504, 16'd3250, 16'd14957, 16'd35521, 16'd32995, 16'd32127, 16'd46679, 16'd18677, 16'd12729}; // indx = 118
    #10;
    addra = 32'd3808;
    dina = {96'd0, 16'd52463, 16'd12269, 16'd21071, 16'd23783, 16'd59414, 16'd30509, 16'd18470, 16'd10789, 16'd13759, 16'd61807}; // indx = 119
    #10;
    addra = 32'd3840;
    dina = {96'd0, 16'd10510, 16'd42412, 16'd57588, 16'd9384, 16'd27356, 16'd27856, 16'd2566, 16'd57662, 16'd31089, 16'd39512}; // indx = 120
    #10;
    addra = 32'd3872;
    dina = {96'd0, 16'd23340, 16'd61589, 16'd43377, 16'd51868, 16'd18524, 16'd23960, 16'd23761, 16'd53109, 16'd8914, 16'd24687}; // indx = 121
    #10;
    addra = 32'd3904;
    dina = {96'd0, 16'd48359, 16'd23888, 16'd20903, 16'd45171, 16'd1778, 16'd14762, 16'd33710, 16'd53871, 16'd13796, 16'd13405}; // indx = 122
    #10;
    addra = 32'd3936;
    dina = {96'd0, 16'd45409, 16'd21362, 16'd13940, 16'd47286, 16'd61062, 16'd54115, 16'd31474, 16'd30933, 16'd16321, 16'd47900}; // indx = 123
    #10;
    addra = 32'd3968;
    dina = {96'd0, 16'd9820, 16'd35320, 16'd6359, 16'd33847, 16'd17743, 16'd10211, 16'd7422, 16'd52251, 16'd18995, 16'd54260}; // indx = 124
    #10;
    addra = 32'd4000;
    dina = {96'd0, 16'd1253, 16'd56388, 16'd56987, 16'd23890, 16'd20052, 16'd16293, 16'd4175, 16'd64339, 16'd17589, 16'd63051}; // indx = 125
    #10;
    addra = 32'd4032;
    dina = {96'd0, 16'd9028, 16'd18208, 16'd60315, 16'd1591, 16'd41189, 16'd61925, 16'd6393, 16'd5543, 16'd43435, 16'd39185}; // indx = 126
    #10;
    addra = 32'd4064;
    dina = {96'd0, 16'd10062, 16'd42477, 16'd12389, 16'd8913, 16'd63896, 16'd31977, 16'd28778, 16'd10595, 16'd39720, 16'd23525}; // indx = 127
    #10;
    addra = 32'd4096;
    dina = {96'd0, 16'd46384, 16'd7992, 16'd55921, 16'd10445, 16'd25170, 16'd43177, 16'd20877, 16'd64022, 16'd6590, 16'd20330}; // indx = 128
    #10;
    addra = 32'd4128;
    dina = {96'd0, 16'd34652, 16'd63844, 16'd48125, 16'd63086, 16'd50368, 16'd52771, 16'd43391, 16'd22813, 16'd7919, 16'd56810}; // indx = 129
    #10;
    addra = 32'd4160;
    dina = {96'd0, 16'd51549, 16'd50228, 16'd62263, 16'd51592, 16'd62894, 16'd3476, 16'd36445, 16'd43646, 16'd41046, 16'd44615}; // indx = 130
    #10;
    addra = 32'd4192;
    dina = {96'd0, 16'd11215, 16'd19246, 16'd45308, 16'd43114, 16'd31923, 16'd62225, 16'd39901, 16'd41263, 16'd46130, 16'd11649}; // indx = 131
    #10;
    addra = 32'd4224;
    dina = {96'd0, 16'd2629, 16'd44031, 16'd7736, 16'd43286, 16'd55381, 16'd18748, 16'd41030, 16'd48593, 16'd10627, 16'd51039}; // indx = 132
    #10;
    addra = 32'd4256;
    dina = {96'd0, 16'd2548, 16'd31115, 16'd19737, 16'd31316, 16'd334, 16'd19758, 16'd17372, 16'd50292, 16'd33511, 16'd34280}; // indx = 133
    #10;
    addra = 32'd4288;
    dina = {96'd0, 16'd36775, 16'd43468, 16'd4112, 16'd19057, 16'd34904, 16'd24480, 16'd53751, 16'd17890, 16'd22822, 16'd26502}; // indx = 134
    #10;
    addra = 32'd4320;
    dina = {96'd0, 16'd4055, 16'd29280, 16'd43690, 16'd24460, 16'd34670, 16'd22910, 16'd52548, 16'd45369, 16'd16869, 16'd3881}; // indx = 135
    #10;
    addra = 32'd4352;
    dina = {96'd0, 16'd48184, 16'd23075, 16'd64569, 16'd32951, 16'd28087, 16'd28085, 16'd55029, 16'd47482, 16'd9388, 16'd30222}; // indx = 136
    #10;
    addra = 32'd4384;
    dina = {96'd0, 16'd23552, 16'd41500, 16'd30784, 16'd1690, 16'd57256, 16'd244, 16'd3120, 16'd11654, 16'd49580, 16'd42369}; // indx = 137
    #10;
    addra = 32'd4416;
    dina = {96'd0, 16'd1160, 16'd6619, 16'd14915, 16'd18416, 16'd31290, 16'd25479, 16'd3047, 16'd4255, 16'd35538, 16'd57189}; // indx = 138
    #10;
    addra = 32'd4448;
    dina = {96'd0, 16'd58707, 16'd47212, 16'd57449, 16'd34945, 16'd16504, 16'd23220, 16'd27638, 16'd36158, 16'd14597, 16'd51187}; // indx = 139
    #10;
    addra = 32'd4480;
    dina = {96'd0, 16'd9088, 16'd62676, 16'd16876, 16'd4191, 16'd23024, 16'd32469, 16'd43094, 16'd55600, 16'd61554, 16'd3855}; // indx = 140
    #10;
    addra = 32'd4512;
    dina = {96'd0, 16'd59007, 16'd51566, 16'd52556, 16'd63700, 16'd31369, 16'd30547, 16'd6346, 16'd45397, 16'd57776, 16'd10115}; // indx = 141
    #10;
    addra = 32'd4544;
    dina = {96'd0, 16'd15700, 16'd14706, 16'd55778, 16'd16012, 16'd47418, 16'd34413, 16'd44035, 16'd16265, 16'd4741, 16'd32754}; // indx = 142
    #10;
    addra = 32'd4576;
    dina = {96'd0, 16'd22308, 16'd372, 16'd60614, 16'd12426, 16'd39015, 16'd56903, 16'd32299, 16'd32839, 16'd40230, 16'd13464}; // indx = 143
    #10;
    addra = 32'd4608;
    dina = {96'd0, 16'd29312, 16'd2093, 16'd10901, 16'd7671, 16'd21846, 16'd9840, 16'd16168, 16'd29670, 16'd41223, 16'd37682}; // indx = 144
    #10;
    addra = 32'd4640;
    dina = {96'd0, 16'd25166, 16'd13838, 16'd44385, 16'd13024, 16'd24395, 16'd5974, 16'd27369, 16'd22927, 16'd46421, 16'd45395}; // indx = 145
    #10;
    addra = 32'd4672;
    dina = {96'd0, 16'd2200, 16'd8535, 16'd65250, 16'd43316, 16'd50701, 16'd20012, 16'd23431, 16'd58241, 16'd18861, 16'd23337}; // indx = 146
    #10;
    addra = 32'd4704;
    dina = {96'd0, 16'd5098, 16'd58545, 16'd21640, 16'd38212, 16'd64949, 16'd53124, 16'd54071, 16'd38217, 16'd41403, 16'd59079}; // indx = 147
    #10;
    addra = 32'd4736;
    dina = {96'd0, 16'd9549, 16'd21671, 16'd42637, 16'd58797, 16'd59177, 16'd48086, 16'd26798, 16'd27605, 16'd51612, 16'd33948}; // indx = 148
    #10;
    addra = 32'd4768;
    dina = {96'd0, 16'd1390, 16'd35082, 16'd56725, 16'd33612, 16'd24286, 16'd27544, 16'd39117, 16'd23407, 16'd64496, 16'd15918}; // indx = 149
    #10;
    addra = 32'd4800;
    dina = {96'd0, 16'd48460, 16'd24846, 16'd18518, 16'd65216, 16'd17547, 16'd7143, 16'd6720, 16'd36513, 16'd16131, 16'd33852}; // indx = 150
    #10;
    addra = 32'd4832;
    dina = {96'd0, 16'd23713, 16'd60687, 16'd30066, 16'd63350, 16'd29892, 16'd29627, 16'd11381, 16'd31905, 16'd60121, 16'd32297}; // indx = 151
    #10;
    addra = 32'd4864;
    dina = {96'd0, 16'd17903, 16'd54104, 16'd56920, 16'd64111, 16'd57779, 16'd30761, 16'd54384, 16'd20491, 16'd329, 16'd4765}; // indx = 152
    #10;
    addra = 32'd4896;
    dina = {96'd0, 16'd28699, 16'd10294, 16'd19165, 16'd2475, 16'd8720, 16'd38308, 16'd345, 16'd28595, 16'd17407, 16'd57228}; // indx = 153
    #10;
    addra = 32'd4928;
    dina = {96'd0, 16'd27945, 16'd37839, 16'd64024, 16'd15969, 16'd52798, 16'd51271, 16'd34257, 16'd40545, 16'd19518, 16'd21331}; // indx = 154
    #10;
    addra = 32'd4960;
    dina = {96'd0, 16'd2862, 16'd15388, 16'd29531, 16'd37486, 16'd64308, 16'd42775, 16'd47392, 16'd38774, 16'd14458, 16'd3408}; // indx = 155
    #10;
    addra = 32'd4992;
    dina = {96'd0, 16'd51367, 16'd43229, 16'd12344, 16'd13952, 16'd4304, 16'd22768, 16'd63564, 16'd17092, 16'd26438, 16'd37709}; // indx = 156
    #10;
    addra = 32'd5024;
    dina = {96'd0, 16'd60857, 16'd63712, 16'd52811, 16'd56061, 16'd5511, 16'd27386, 16'd18911, 16'd61954, 16'd59946, 16'd18501}; // indx = 157
    #10;
    addra = 32'd5056;
    dina = {96'd0, 16'd48368, 16'd25146, 16'd13852, 16'd12246, 16'd64825, 16'd18564, 16'd16253, 16'd61315, 16'd50544, 16'd26106}; // indx = 158
    #10;
    addra = 32'd5088;
    dina = {96'd0, 16'd8118, 16'd24357, 16'd3413, 16'd16578, 16'd10563, 16'd57860, 16'd1041, 16'd32588, 16'd39197, 16'd12851}; // indx = 159
    #10;
    addra = 32'd5120;
    dina = {96'd0, 16'd57286, 16'd61824, 16'd51158, 16'd45247, 16'd62121, 16'd17593, 16'd59940, 16'd11416, 16'd28006, 16'd15959}; // indx = 160
    #10;
    addra = 32'd5152;
    dina = {96'd0, 16'd17774, 16'd19507, 16'd12460, 16'd22998, 16'd9074, 16'd42450, 16'd16118, 16'd12013, 16'd20743, 16'd40730}; // indx = 161
    #10;
    addra = 32'd5184;
    dina = {96'd0, 16'd32459, 16'd4843, 16'd2442, 16'd56512, 16'd29831, 16'd3490, 16'd7048, 16'd25159, 16'd10357, 16'd25131}; // indx = 162
    #10;
    addra = 32'd5216;
    dina = {96'd0, 16'd50487, 16'd5397, 16'd63373, 16'd45438, 16'd50192, 16'd24747, 16'd39081, 16'd54855, 16'd25577, 16'd65106}; // indx = 163
    #10;
    addra = 32'd5248;
    dina = {96'd0, 16'd9840, 16'd25068, 16'd30637, 16'd61932, 16'd49839, 16'd48029, 16'd51650, 16'd34601, 16'd57191, 16'd5779}; // indx = 164
    #10;
    addra = 32'd5280;
    dina = {96'd0, 16'd34061, 16'd47094, 16'd28974, 16'd64395, 16'd58006, 16'd51147, 16'd46188, 16'd41654, 16'd59272, 16'd42866}; // indx = 165
    #10;
    addra = 32'd5312;
    dina = {96'd0, 16'd15887, 16'd49965, 16'd35019, 16'd30597, 16'd64107, 16'd17797, 16'd47073, 16'd12462, 16'd31789, 16'd7916}; // indx = 166
    #10;
    addra = 32'd5344;
    dina = {96'd0, 16'd42394, 16'd25580, 16'd30721, 16'd54086, 16'd28571, 16'd54955, 16'd28045, 16'd44763, 16'd47241, 16'd7225}; // indx = 167
    #10;
    addra = 32'd5376;
    dina = {96'd0, 16'd65373, 16'd44537, 16'd36288, 16'd59500, 16'd48598, 16'd12879, 16'd53547, 16'd61083, 16'd38877, 16'd3264}; // indx = 168
    #10;
    addra = 32'd5408;
    dina = {96'd0, 16'd27367, 16'd49810, 16'd60525, 16'd18976, 16'd24401, 16'd25455, 16'd5904, 16'd22393, 16'd42040, 16'd48529}; // indx = 169
    #10;
    addra = 32'd5440;
    dina = {96'd0, 16'd60858, 16'd27382, 16'd54658, 16'd2123, 16'd39358, 16'd11849, 16'd38432, 16'd42838, 16'd55400, 16'd62263}; // indx = 170
    #10;
    addra = 32'd5472;
    dina = {96'd0, 16'd2484, 16'd3624, 16'd22821, 16'd61013, 16'd18361, 16'd25604, 16'd7289, 16'd58457, 16'd9256, 16'd50942}; // indx = 171
    #10;
    addra = 32'd5504;
    dina = {96'd0, 16'd12012, 16'd48484, 16'd44453, 16'd34523, 16'd57685, 16'd3444, 16'd2817, 16'd35777, 16'd31498, 16'd57245}; // indx = 172
    #10;
    addra = 32'd5536;
    dina = {96'd0, 16'd30658, 16'd37802, 16'd11742, 16'd40104, 16'd19929, 16'd36312, 16'd50528, 16'd57760, 16'd51118, 16'd65262}; // indx = 173
    #10;
    addra = 32'd5568;
    dina = {96'd0, 16'd32922, 16'd5865, 16'd34775, 16'd46965, 16'd18441, 16'd62210, 16'd41702, 16'd53169, 16'd46281, 16'd6364}; // indx = 174
    #10;
    addra = 32'd5600;
    dina = {96'd0, 16'd62275, 16'd21735, 16'd28325, 16'd17764, 16'd11229, 16'd45288, 16'd15594, 16'd26710, 16'd25632, 16'd6714}; // indx = 175
    #10;
    addra = 32'd5632;
    dina = {96'd0, 16'd27037, 16'd57551, 16'd37465, 16'd37168, 16'd3417, 16'd60523, 16'd20323, 16'd3638, 16'd60700, 16'd58180}; // indx = 176
    #10;
    addra = 32'd5664;
    dina = {96'd0, 16'd1312, 16'd54448, 16'd13204, 16'd32216, 16'd63214, 16'd10536, 16'd37666, 16'd27999, 16'd51211, 16'd14967}; // indx = 177
    #10;
    addra = 32'd5696;
    dina = {96'd0, 16'd52495, 16'd26090, 16'd63925, 16'd19490, 16'd53735, 16'd16794, 16'd15171, 16'd16785, 16'd50381, 16'd24940}; // indx = 178
    #10;
    addra = 32'd5728;
    dina = {96'd0, 16'd8375, 16'd63977, 16'd64072, 16'd41362, 16'd22870, 16'd24091, 16'd36601, 16'd8157, 16'd57811, 16'd34203}; // indx = 179
    #10;
    addra = 32'd5760;
    dina = {96'd0, 16'd60166, 16'd2575, 16'd41679, 16'd7189, 16'd29249, 16'd31364, 16'd47389, 16'd2464, 16'd12714, 16'd25463}; // indx = 180
    #10;
    addra = 32'd5792;
    dina = {96'd0, 16'd52278, 16'd16062, 16'd62490, 16'd46732, 16'd46216, 16'd37927, 16'd17844, 16'd54276, 16'd55423, 16'd2732}; // indx = 181
    #10;
    addra = 32'd5824;
    dina = {96'd0, 16'd44767, 16'd62734, 16'd43324, 16'd28513, 16'd16710, 16'd45550, 16'd18255, 16'd57144, 16'd2905, 16'd43666}; // indx = 182
    #10;
    addra = 32'd5856;
    dina = {96'd0, 16'd65277, 16'd63979, 16'd18854, 16'd12713, 16'd42282, 16'd59069, 16'd48669, 16'd60991, 16'd6298, 16'd31540}; // indx = 183
    #10;
    addra = 32'd5888;
    dina = {96'd0, 16'd7827, 16'd10019, 16'd48750, 16'd10818, 16'd6900, 16'd63402, 16'd51483, 16'd43933, 16'd24179, 16'd9440}; // indx = 184
    #10;
    addra = 32'd5920;
    dina = {96'd0, 16'd61962, 16'd806, 16'd63792, 16'd30713, 16'd35646, 16'd26738, 16'd33127, 16'd41262, 16'd54140, 16'd39242}; // indx = 185
    #10;
    addra = 32'd5952;
    dina = {96'd0, 16'd41514, 16'd11812, 16'd9563, 16'd21064, 16'd53421, 16'd50056, 16'd22033, 16'd47536, 16'd23768, 16'd55339}; // indx = 186
    #10;
    addra = 32'd5984;
    dina = {96'd0, 16'd33320, 16'd26537, 16'd58631, 16'd47279, 16'd59868, 16'd34484, 16'd62626, 16'd10227, 16'd23491, 16'd60735}; // indx = 187
    #10;
    addra = 32'd6016;
    dina = {96'd0, 16'd9613, 16'd24298, 16'd48898, 16'd32810, 16'd34341, 16'd44801, 16'd61714, 16'd7177, 16'd29630, 16'd21783}; // indx = 188
    #10;
    addra = 32'd6048;
    dina = {96'd0, 16'd52628, 16'd22099, 16'd44595, 16'd18023, 16'd13607, 16'd51149, 16'd7282, 16'd61611, 16'd40458, 16'd16197}; // indx = 189
    #10;
    addra = 32'd6080;
    dina = {96'd0, 16'd5035, 16'd26372, 16'd10159, 16'd22219, 16'd10196, 16'd52570, 16'd50625, 16'd26485, 16'd60314, 16'd57813}; // indx = 190
    #10;
    addra = 32'd6112;
    dina = {96'd0, 16'd38670, 16'd47985, 16'd55819, 16'd22142, 16'd49996, 16'd58244, 16'd44214, 16'd39058, 16'd394, 16'd11083}; // indx = 191
    #10;
    addra = 32'd6144;
    dina = {96'd0, 16'd524, 16'd578, 16'd58300, 16'd1949, 16'd59308, 16'd46992, 16'd30222, 16'd10369, 16'd34102, 16'd41826}; // indx = 192
    #10;
    addra = 32'd6176;
    dina = {96'd0, 16'd42530, 16'd27103, 16'd15711, 16'd64626, 16'd59397, 16'd1319, 16'd12645, 16'd252, 16'd21002, 16'd38009}; // indx = 193
    #10;
    addra = 32'd6208;
    dina = {96'd0, 16'd2617, 16'd21125, 16'd24348, 16'd24021, 16'd35065, 16'd27340, 16'd34628, 16'd15017, 16'd34071, 16'd64585}; // indx = 194
    #10;
    addra = 32'd6240;
    dina = {96'd0, 16'd55534, 16'd62097, 16'd58591, 16'd62871, 16'd48576, 16'd45610, 16'd26918, 16'd62882, 16'd41833, 16'd3223}; // indx = 195
    #10;
    addra = 32'd6272;
    dina = {96'd0, 16'd41853, 16'd19459, 16'd45478, 16'd23349, 16'd45468, 16'd63972, 16'd33318, 16'd33820, 16'd47448, 16'd58126}; // indx = 196
    #10;
    addra = 32'd6304;
    dina = {96'd0, 16'd49863, 16'd37909, 16'd27623, 16'd42196, 16'd34930, 16'd13166, 16'd56408, 16'd21909, 16'd37410, 16'd1306}; // indx = 197
    #10;
    addra = 32'd6336;
    dina = {96'd0, 16'd17710, 16'd45527, 16'd4708, 16'd16032, 16'd5511, 16'd34657, 16'd1558, 16'd1110, 16'd51286, 16'd48265}; // indx = 198
    #10;
    addra = 32'd6368;
    dina = {96'd0, 16'd56573, 16'd4743, 16'd24956, 16'd16734, 16'd7715, 16'd22829, 16'd35837, 16'd54362, 16'd10169, 16'd63243}; // indx = 199
    #10;
    addra = 32'd6400;
    dina = {96'd0, 16'd43636, 16'd60531, 16'd45176, 16'd8041, 16'd6531, 16'd50083, 16'd5789, 16'd42737, 16'd57192, 16'd50725}; // indx = 200
    #10;
    addra = 32'd6432;
    dina = {96'd0, 16'd56200, 16'd27042, 16'd36841, 16'd44190, 16'd25859, 16'd12150, 16'd5590, 16'd19605, 16'd32807, 16'd16260}; // indx = 201
    #10;
    addra = 32'd6464;
    dina = {96'd0, 16'd63632, 16'd24268, 16'd47792, 16'd1577, 16'd60304, 16'd12945, 16'd12960, 16'd60921, 16'd63700, 16'd53070}; // indx = 202
    #10;
    addra = 32'd6496;
    dina = {96'd0, 16'd8428, 16'd42488, 16'd13306, 16'd46081, 16'd33856, 16'd61159, 16'd23406, 16'd15918, 16'd12548, 16'd64992}; // indx = 203
    #10;
    addra = 32'd6528;
    dina = {96'd0, 16'd48404, 16'd38285, 16'd24600, 16'd42050, 16'd43479, 16'd875, 16'd25770, 16'd58483, 16'd25802, 16'd6439}; // indx = 204
    #10;
    addra = 32'd6560;
    dina = {96'd0, 16'd12732, 16'd54772, 16'd9720, 16'd18207, 16'd18765, 16'd55253, 16'd49665, 16'd22868, 16'd42204, 16'd62818}; // indx = 205
    #10;
    addra = 32'd6592;
    dina = {96'd0, 16'd44108, 16'd50479, 16'd38712, 16'd49094, 16'd40804, 16'd33238, 16'd59329, 16'd25825, 16'd6323, 16'd1594}; // indx = 206
    #10;
    addra = 32'd6624;
    dina = {96'd0, 16'd14668, 16'd7768, 16'd61712, 16'd14528, 16'd6442, 16'd54252, 16'd53154, 16'd24408, 16'd50326, 16'd6923}; // indx = 207
    #10;
    addra = 32'd6656;
    dina = {96'd0, 16'd60599, 16'd10049, 16'd19619, 16'd20683, 16'd54844, 16'd2486, 16'd49541, 16'd39019, 16'd30627, 16'd3101}; // indx = 208
    #10;
    addra = 32'd6688;
    dina = {96'd0, 16'd17120, 16'd2162, 16'd34995, 16'd4762, 16'd61900, 16'd63833, 16'd33542, 16'd34866, 16'd33922, 16'd61705}; // indx = 209
    #10;
    addra = 32'd6720;
    dina = {96'd0, 16'd13984, 16'd4336, 16'd57490, 16'd22313, 16'd52254, 16'd21078, 16'd17439, 16'd8959, 16'd13395, 16'd51312}; // indx = 210
    #10;
    addra = 32'd6752;
    dina = {96'd0, 16'd10003, 16'd35525, 16'd57623, 16'd3726, 16'd56616, 16'd55435, 16'd50509, 16'd46785, 16'd24241, 16'd43246}; // indx = 211
    #10;
    addra = 32'd6784;
    dina = {96'd0, 16'd48874, 16'd17801, 16'd43287, 16'd4747, 16'd16990, 16'd37439, 16'd3374, 16'd26590, 16'd39928, 16'd36734}; // indx = 212
    #10;
    addra = 32'd6816;
    dina = {96'd0, 16'd26047, 16'd15947, 16'd24747, 16'd25206, 16'd18747, 16'd57455, 16'd33375, 16'd33629, 16'd7373, 16'd40090}; // indx = 213
    #10;
    addra = 32'd6848;
    dina = {96'd0, 16'd28776, 16'd1985, 16'd64140, 16'd24323, 16'd4359, 16'd525, 16'd53884, 16'd6084, 16'd17784, 16'd35306}; // indx = 214
    #10;
    addra = 32'd6880;
    dina = {96'd0, 16'd32048, 16'd11864, 16'd27215, 16'd54815, 16'd23685, 16'd55647, 16'd31084, 16'd4432, 16'd55949, 16'd26027}; // indx = 215
    #10;
    addra = 32'd6912;
    dina = {96'd0, 16'd49568, 16'd9190, 16'd38665, 16'd21017, 16'd11361, 16'd13566, 16'd43157, 16'd949, 16'd51434, 16'd16845}; // indx = 216
    #10;
    addra = 32'd6944;
    dina = {96'd0, 16'd47537, 16'd63152, 16'd55659, 16'd49431, 16'd10144, 16'd54053, 16'd4920, 16'd44111, 16'd8966, 16'd36911}; // indx = 217
    #10;
    addra = 32'd6976;
    dina = {96'd0, 16'd38710, 16'd21259, 16'd9702, 16'd34573, 16'd48269, 16'd7660, 16'd41238, 16'd48672, 16'd19508, 16'd17484}; // indx = 218
    #10;
    addra = 32'd7008;
    dina = {96'd0, 16'd31682, 16'd58478, 16'd46865, 16'd46913, 16'd49952, 16'd53780, 16'd45617, 16'd40467, 16'd42814, 16'd2930}; // indx = 219
    #10;
    addra = 32'd7040;
    dina = {96'd0, 16'd55928, 16'd64920, 16'd15757, 16'd36528, 16'd1875, 16'd29952, 16'd3694, 16'd64100, 16'd49385, 16'd31995}; // indx = 220
    #10;
    addra = 32'd7072;
    dina = {96'd0, 16'd23046, 16'd23785, 16'd28096, 16'd29117, 16'd33080, 16'd8302, 16'd31906, 16'd62639, 16'd32367, 16'd49310}; // indx = 221
    #10;
    addra = 32'd7104;
    dina = {96'd0, 16'd14375, 16'd19009, 16'd27377, 16'd46478, 16'd32793, 16'd7346, 16'd65191, 16'd34529, 16'd47192, 16'd3065}; // indx = 222
    #10;
    addra = 32'd7136;
    dina = {96'd0, 16'd34464, 16'd45683, 16'd34997, 16'd52154, 16'd57987, 16'd51519, 16'd39846, 16'd58229, 16'd2124, 16'd12513}; // indx = 223
    #10;
    addra = 32'd7168;
    dina = {96'd0, 16'd6285, 16'd26806, 16'd55477, 16'd16833, 16'd15997, 16'd15921, 16'd65178, 16'd28282, 16'd58762, 16'd13173}; // indx = 224
    #10;
    addra = 32'd7200;
    dina = {96'd0, 16'd32894, 16'd54799, 16'd59841, 16'd2624, 16'd37611, 16'd14024, 16'd33619, 16'd57577, 16'd3048, 16'd63127}; // indx = 225
    #10;
    addra = 32'd7232;
    dina = {96'd0, 16'd64194, 16'd18574, 16'd3719, 16'd27810, 16'd22907, 16'd30991, 16'd36030, 16'd17623, 16'd26979, 16'd12451}; // indx = 226
    #10;
    addra = 32'd7264;
    dina = {96'd0, 16'd37852, 16'd23271, 16'd5393, 16'd15303, 16'd21852, 16'd62087, 16'd16018, 16'd14993, 16'd45460, 16'd57982}; // indx = 227
    #10;
    addra = 32'd7296;
    dina = {96'd0, 16'd12277, 16'd14617, 16'd60364, 16'd25797, 16'd61822, 16'd13911, 16'd45948, 16'd3697, 16'd22565, 16'd14189}; // indx = 228
    #10;
    addra = 32'd7328;
    dina = {96'd0, 16'd5074, 16'd5603, 16'd19713, 16'd21814, 16'd61352, 16'd56511, 16'd15993, 16'd26339, 16'd61740, 16'd9580}; // indx = 229
    #10;
    addra = 32'd7360;
    dina = {96'd0, 16'd36009, 16'd59273, 16'd16728, 16'd35776, 16'd32898, 16'd63520, 16'd60801, 16'd39211, 16'd28821, 16'd12160}; // indx = 230
    #10;
    addra = 32'd7392;
    dina = {96'd0, 16'd51361, 16'd15075, 16'd54833, 16'd57104, 16'd31027, 16'd24409, 16'd5617, 16'd22728, 16'd52963, 16'd64798}; // indx = 231
    #10;
    addra = 32'd7424;
    dina = {96'd0, 16'd25937, 16'd54797, 16'd59463, 16'd52758, 16'd24978, 16'd39972, 16'd32645, 16'd27681, 16'd58280, 16'd14489}; // indx = 232
    #10;
    addra = 32'd7456;
    dina = {96'd0, 16'd6765, 16'd11191, 16'd52558, 16'd54010, 16'd53352, 16'd30565, 16'd48452, 16'd32095, 16'd21030, 16'd50845}; // indx = 233
    #10;
    addra = 32'd7488;
    dina = {96'd0, 16'd28932, 16'd22560, 16'd55008, 16'd36915, 16'd16352, 16'd25108, 16'd6810, 16'd51997, 16'd24025, 16'd62944}; // indx = 234
    #10;
    addra = 32'd7520;
    dina = {96'd0, 16'd12732, 16'd25297, 16'd30605, 16'd35618, 16'd23132, 16'd48639, 16'd38340, 16'd25429, 16'd38258, 16'd46496}; // indx = 235
    #10;
    addra = 32'd7552;
    dina = {96'd0, 16'd5710, 16'd4132, 16'd50892, 16'd10722, 16'd2334, 16'd41113, 16'd23008, 16'd53814, 16'd36884, 16'd24715}; // indx = 236
    #10;
    addra = 32'd7584;
    dina = {96'd0, 16'd65385, 16'd58191, 16'd45253, 16'd50395, 16'd25306, 16'd59540, 16'd38885, 16'd61684, 16'd64801, 16'd32613}; // indx = 237
    #10;
    addra = 32'd7616;
    dina = {96'd0, 16'd14396, 16'd12742, 16'd46123, 16'd35104, 16'd47649, 16'd3941, 16'd83, 16'd5696, 16'd48467, 16'd31845}; // indx = 238
    #10;
    addra = 32'd7648;
    dina = {96'd0, 16'd29042, 16'd59063, 16'd3515, 16'd47351, 16'd59646, 16'd26821, 16'd20902, 16'd60194, 16'd60830, 16'd41302}; // indx = 239
    #10;
    addra = 32'd7680;
    dina = {96'd0, 16'd60422, 16'd34600, 16'd10062, 16'd10033, 16'd45271, 16'd33848, 16'd23315, 16'd8781, 16'd1588, 16'd56155}; // indx = 240
    #10;
    addra = 32'd7712;
    dina = {96'd0, 16'd31521, 16'd20676, 16'd21150, 16'd16987, 16'd19151, 16'd52308, 16'd26776, 16'd47043, 16'd2559, 16'd16909}; // indx = 241
    #10;
    addra = 32'd7744;
    dina = {96'd0, 16'd4018, 16'd8110, 16'd42165, 16'd9764, 16'd6735, 16'd48133, 16'd4450, 16'd59553, 16'd28507, 16'd51008}; // indx = 242
    #10;
    addra = 32'd7776;
    dina = {96'd0, 16'd50373, 16'd63535, 16'd29755, 16'd64771, 16'd39652, 16'd14716, 16'd47518, 16'd23657, 16'd59684, 16'd18183}; // indx = 243
    #10;
    addra = 32'd7808;
    dina = {96'd0, 16'd4848, 16'd34570, 16'd40740, 16'd59469, 16'd14208, 16'd16585, 16'd19420, 16'd31563, 16'd6356, 16'd27862}; // indx = 244
    #10;
    addra = 32'd7840;
    dina = {96'd0, 16'd56382, 16'd65144, 16'd911, 16'd51057, 16'd56275, 16'd5785, 16'd11343, 16'd7535, 16'd55810, 16'd21523}; // indx = 245
    #10;
    addra = 32'd7872;
    dina = {96'd0, 16'd15034, 16'd9967, 16'd36129, 16'd24363, 16'd17916, 16'd49331, 16'd62133, 16'd58633, 16'd36098, 16'd52601}; // indx = 246
    #10;
    addra = 32'd7904;
    dina = {96'd0, 16'd64694, 16'd39336, 16'd19426, 16'd26888, 16'd54260, 16'd29525, 16'd47058, 16'd18312, 16'd32497, 16'd62568}; // indx = 247
    #10;
    addra = 32'd7936;
    dina = {96'd0, 16'd60390, 16'd63062, 16'd13472, 16'd42077, 16'd24777, 16'd48873, 16'd13526, 16'd28643, 16'd12701, 16'd26124}; // indx = 248
    #10;
    addra = 32'd7968;
    dina = {96'd0, 16'd11563, 16'd2847, 16'd43161, 16'd9374, 16'd62467, 16'd5050, 16'd21093, 16'd12120, 16'd13640, 16'd2361}; // indx = 249
    #10;
    addra = 32'd8000;
    dina = {96'd0, 16'd52211, 16'd52612, 16'd65460, 16'd47860, 16'd27981, 16'd54064, 16'd419, 16'd9140, 16'd58174, 16'd38112}; // indx = 250
    #10;
    addra = 32'd8032;
    dina = {96'd0, 16'd38595, 16'd18455, 16'd58295, 16'd63484, 16'd24874, 16'd63134, 16'd55178, 16'd23277, 16'd54666, 16'd15751}; // indx = 251
    #10;
    addra = 32'd8064;
    dina = {96'd0, 16'd13268, 16'd19283, 16'd38543, 16'd51371, 16'd57514, 16'd29090, 16'd6764, 16'd47317, 16'd37094, 16'd42022}; // indx = 252
    #10;
    addra = 32'd8096;
    dina = {96'd0, 16'd49923, 16'd9023, 16'd37475, 16'd8942, 16'd23405, 16'd36043, 16'd6248, 16'd28159, 16'd46215, 16'd50009}; // indx = 253
    #10;
    addra = 32'd8128;
    dina = {96'd0, 16'd28265, 16'd53719, 16'd37676, 16'd21752, 16'd6480, 16'd1029, 16'd3142, 16'd35483, 16'd11636, 16'd20637}; // indx = 254
    #10;
    addra = 32'd8160;
    dina = {96'd0, 16'd39492, 16'd48558, 16'd56348, 16'd13985, 16'd54532, 16'd59362, 16'd47745, 16'd31644, 16'd36071, 16'd49231}; // indx = 255
    #10;
    addra = 32'd8192;
    dina = {96'd0, 16'd29319, 16'd29712, 16'd65051, 16'd64762, 16'd22565, 16'd36350, 16'd64118, 16'd16153, 16'd64885, 16'd12946}; // indx = 256
    #10;
    addra = 32'd8224;
    dina = {96'd0, 16'd6531, 16'd36299, 16'd18461, 16'd9442, 16'd60188, 16'd62389, 16'd53836, 16'd44496, 16'd46382, 16'd31475}; // indx = 257
    #10;
    addra = 32'd8256;
    dina = {96'd0, 16'd53080, 16'd62425, 16'd57678, 16'd55006, 16'd21581, 16'd12176, 16'd60289, 16'd15218, 16'd52908, 16'd16843}; // indx = 258
    #10;
    addra = 32'd8288;
    dina = {96'd0, 16'd17113, 16'd15931, 16'd65402, 16'd19270, 16'd10725, 16'd34156, 16'd57759, 16'd43198, 16'd42605, 16'd15845}; // indx = 259
    #10;
    addra = 32'd8320;
    dina = {96'd0, 16'd2860, 16'd9834, 16'd50214, 16'd6457, 16'd18020, 16'd2974, 16'd58708, 16'd14756, 16'd41860, 16'd16677}; // indx = 260
    #10;
    addra = 32'd8352;
    dina = {96'd0, 16'd43035, 16'd13397, 16'd46062, 16'd303, 16'd61778, 16'd6125, 16'd35533, 16'd29570, 16'd21426, 16'd46230}; // indx = 261
    #10;
    addra = 32'd8384;
    dina = {96'd0, 16'd10521, 16'd22848, 16'd12700, 16'd15902, 16'd12329, 16'd63870, 16'd61191, 16'd59229, 16'd53434, 16'd46161}; // indx = 262
    #10;
    addra = 32'd8416;
    dina = {96'd0, 16'd58392, 16'd9597, 16'd41229, 16'd45633, 16'd26290, 16'd50674, 16'd51623, 16'd17154, 16'd56841, 16'd19023}; // indx = 263
    #10;
    addra = 32'd8448;
    dina = {96'd0, 16'd51833, 16'd25116, 16'd39195, 16'd63826, 16'd15570, 16'd18033, 16'd48120, 16'd51992, 16'd21090, 16'd27236}; // indx = 264
    #10;
    addra = 32'd8480;
    dina = {96'd0, 16'd17633, 16'd12418, 16'd35489, 16'd62389, 16'd54123, 16'd50027, 16'd61903, 16'd12514, 16'd16608, 16'd30587}; // indx = 265
    #10;
    addra = 32'd8512;
    dina = {96'd0, 16'd59564, 16'd51323, 16'd62876, 16'd40558, 16'd61587, 16'd62529, 16'd37237, 16'd54239, 16'd39800, 16'd44790}; // indx = 266
    #10;
    addra = 32'd8544;
    dina = {96'd0, 16'd13788, 16'd64186, 16'd26521, 16'd64199, 16'd7461, 16'd43339, 16'd21042, 16'd54452, 16'd52662, 16'd12998}; // indx = 267
    #10;
    addra = 32'd8576;
    dina = {96'd0, 16'd36451, 16'd26468, 16'd38674, 16'd54179, 16'd3233, 16'd59493, 16'd47697, 16'd32492, 16'd11586, 16'd41711}; // indx = 268
    #10;
    addra = 32'd8608;
    dina = {96'd0, 16'd49642, 16'd51142, 16'd52712, 16'd6015, 16'd4688, 16'd13889, 16'd22733, 16'd53467, 16'd64264, 16'd14089}; // indx = 269
    #10;
    addra = 32'd8640;
    dina = {96'd0, 16'd8165, 16'd31132, 16'd42658, 16'd17232, 16'd21748, 16'd62093, 16'd56090, 16'd27788, 16'd52932, 16'd24468}; // indx = 270
    #10;
    addra = 32'd8672;
    dina = {96'd0, 16'd34847, 16'd29030, 16'd9909, 16'd5562, 16'd5751, 16'd52370, 16'd57698, 16'd30719, 16'd10862, 16'd6335}; // indx = 271
    #10;
    addra = 32'd8704;
    dina = {96'd0, 16'd45662, 16'd51950, 16'd35058, 16'd24293, 16'd14029, 16'd56022, 16'd4996, 16'd43384, 16'd14566, 16'd38347}; // indx = 272
    #10;
    addra = 32'd8736;
    dina = {96'd0, 16'd544, 16'd40583, 16'd21228, 16'd27052, 16'd1479, 16'd43567, 16'd4418, 16'd26923, 16'd40435, 16'd25255}; // indx = 273
    #10;
    addra = 32'd8768;
    dina = {96'd0, 16'd15447, 16'd39935, 16'd7775, 16'd29210, 16'd25204, 16'd43713, 16'd13976, 16'd53784, 16'd54419, 16'd53860}; // indx = 274
    #10;
    addra = 32'd8800;
    dina = {96'd0, 16'd12274, 16'd51910, 16'd39902, 16'd9783, 16'd41068, 16'd6263, 16'd57564, 16'd5677, 16'd59180, 16'd35890}; // indx = 275
    #10;
    addra = 32'd8832;
    dina = {96'd0, 16'd10047, 16'd4424, 16'd52266, 16'd61420, 16'd49197, 16'd52267, 16'd37916, 16'd27797, 16'd59732, 16'd31896}; // indx = 276
    #10;
    addra = 32'd8864;
    dina = {96'd0, 16'd7378, 16'd40415, 16'd35330, 16'd6657, 16'd10243, 16'd31399, 16'd23892, 16'd18789, 16'd58716, 16'd39947}; // indx = 277
    #10;
    addra = 32'd8896;
    dina = {96'd0, 16'd8708, 16'd582, 16'd11872, 16'd26085, 16'd52336, 16'd17782, 16'd40573, 16'd23623, 16'd22401, 16'd25457}; // indx = 278
    #10;
    addra = 32'd8928;
    dina = {96'd0, 16'd47908, 16'd4046, 16'd39766, 16'd2576, 16'd14464, 16'd17932, 16'd62204, 16'd12493, 16'd1029, 16'd40082}; // indx = 279
    #10;
    addra = 32'd8960;
    dina = {96'd0, 16'd53895, 16'd31252, 16'd11202, 16'd20699, 16'd65380, 16'd42059, 16'd42731, 16'd48678, 16'd11752, 16'd36801}; // indx = 280
    #10;
    addra = 32'd8992;
    dina = {96'd0, 16'd4770, 16'd28497, 16'd21900, 16'd28875, 16'd62648, 16'd15154, 16'd55114, 16'd5167, 16'd12307, 16'd4143}; // indx = 281
    #10;
    addra = 32'd9024;
    dina = {96'd0, 16'd45425, 16'd43811, 16'd39533, 16'd663, 16'd10522, 16'd10629, 16'd30138, 16'd1059, 16'd20211, 16'd23487}; // indx = 282
    #10;
    addra = 32'd9056;
    dina = {96'd0, 16'd7573, 16'd42098, 16'd13009, 16'd31554, 16'd45824, 16'd34522, 16'd16008, 16'd44486, 16'd44425, 16'd38845}; // indx = 283
    #10;
    addra = 32'd9088;
    dina = {96'd0, 16'd23371, 16'd44659, 16'd24118, 16'd29938, 16'd27330, 16'd36048, 16'd60937, 16'd8939, 16'd54669, 16'd12024}; // indx = 284
    #10;
    addra = 32'd9120;
    dina = {96'd0, 16'd13033, 16'd10494, 16'd40056, 16'd7895, 16'd26119, 16'd1224, 16'd7403, 16'd46313, 16'd63671, 16'd28506}; // indx = 285
    #10;
    addra = 32'd9152;
    dina = {96'd0, 16'd13412, 16'd30558, 16'd53668, 16'd31770, 16'd12097, 16'd15070, 16'd25871, 16'd58059, 16'd63243, 16'd11100}; // indx = 286
    #10;
    addra = 32'd9184;
    dina = {96'd0, 16'd36240, 16'd43541, 16'd45903, 16'd37382, 16'd24602, 16'd31122, 16'd351, 16'd38024, 16'd31527, 16'd21863}; // indx = 287
    #10;
    addra = 32'd9216;
    dina = {96'd0, 16'd46528, 16'd39138, 16'd9400, 16'd62241, 16'd2688, 16'd22760, 16'd4441, 16'd64108, 16'd51394, 16'd23726}; // indx = 288
    #10;
    addra = 32'd9248;
    dina = {96'd0, 16'd50630, 16'd36658, 16'd65141, 16'd29261, 16'd3695, 16'd1500, 16'd4927, 16'd7162, 16'd50559, 16'd14073}; // indx = 289
    #10;
    addra = 32'd9280;
    dina = {96'd0, 16'd7552, 16'd45287, 16'd17376, 16'd55438, 16'd31336, 16'd56572, 16'd4582, 16'd3550, 16'd60087, 16'd53742}; // indx = 290
    #10;
    addra = 32'd9312;
    dina = {96'd0, 16'd52251, 16'd9591, 16'd53192, 16'd31067, 16'd57579, 16'd5705, 16'd21923, 16'd28642, 16'd46612, 16'd767}; // indx = 291
    #10;
    addra = 32'd9344;
    dina = {96'd0, 16'd15978, 16'd30327, 16'd44135, 16'd10502, 16'd19229, 16'd11057, 16'd46854, 16'd48714, 16'd64861, 16'd19692}; // indx = 292
    #10;
    addra = 32'd9376;
    dina = {96'd0, 16'd14449, 16'd5082, 16'd28481, 16'd56439, 16'd29721, 16'd8777, 16'd39261, 16'd64831, 16'd33972, 16'd20640}; // indx = 293
    #10;
    addra = 32'd9408;
    dina = {96'd0, 16'd17832, 16'd62090, 16'd21137, 16'd44639, 16'd30542, 16'd23006, 16'd10104, 16'd44662, 16'd52879, 16'd43009}; // indx = 294
    #10;
    addra = 32'd9440;
    dina = {96'd0, 16'd52581, 16'd23571, 16'd19157, 16'd45596, 16'd13496, 16'd4383, 16'd6744, 16'd31014, 16'd12370, 16'd40024}; // indx = 295
    #10;
    addra = 32'd9472;
    dina = {96'd0, 16'd58325, 16'd17245, 16'd27110, 16'd54352, 16'd117, 16'd42164, 16'd9113, 16'd41827, 16'd17114, 16'd25971}; // indx = 296
    #10;
    addra = 32'd9504;
    dina = {96'd0, 16'd1625, 16'd58798, 16'd10573, 16'd64471, 16'd38006, 16'd48911, 16'd59974, 16'd54831, 16'd51961, 16'd20980}; // indx = 297
    #10;
    addra = 32'd9536;
    dina = {96'd0, 16'd35465, 16'd54323, 16'd37205, 16'd46574, 16'd63901, 16'd22646, 16'd25457, 16'd41329, 16'd25221, 16'd18851}; // indx = 298
    #10;
    addra = 32'd9568;
    dina = {96'd0, 16'd46461, 16'd13969, 16'd58860, 16'd37743, 16'd14478, 16'd344, 16'd41509, 16'd52427, 16'd43111, 16'd19377}; // indx = 299
    #10;
    addra = 32'd9600;
    dina = {96'd0, 16'd53363, 16'd39348, 16'd21890, 16'd6618, 16'd45831, 16'd7169, 16'd451, 16'd3945, 16'd56907, 16'd63965}; // indx = 300
    #10;
    addra = 32'd9632;
    dina = {96'd0, 16'd49360, 16'd48914, 16'd45743, 16'd5932, 16'd11677, 16'd56642, 16'd22558, 16'd11395, 16'd22275, 16'd45154}; // indx = 301
    #10;
    addra = 32'd9664;
    dina = {96'd0, 16'd45258, 16'd16375, 16'd15057, 16'd11061, 16'd54574, 16'd61218, 16'd26912, 16'd61755, 16'd19791, 16'd56495}; // indx = 302
    #10;
    addra = 32'd9696;
    dina = {96'd0, 16'd55959, 16'd12806, 16'd36397, 16'd29665, 16'd32689, 16'd16838, 16'd53835, 16'd19370, 16'd19569, 16'd33838}; // indx = 303
    #10;
    addra = 32'd9728;
    dina = {96'd0, 16'd45572, 16'd2427, 16'd45024, 16'd45236, 16'd6463, 16'd39441, 16'd37219, 16'd32672, 16'd19104, 16'd10228}; // indx = 304
    #10;
    addra = 32'd9760;
    dina = {96'd0, 16'd41928, 16'd12314, 16'd53359, 16'd10675, 16'd20609, 16'd64475, 16'd36218, 16'd12431, 16'd44964, 16'd19569}; // indx = 305
    #10;
    addra = 32'd9792;
    dina = {96'd0, 16'd24283, 16'd21894, 16'd50394, 16'd27186, 16'd51438, 16'd45163, 16'd36350, 16'd10701, 16'd53663, 16'd5567}; // indx = 306
    #10;
    addra = 32'd9824;
    dina = {96'd0, 16'd51724, 16'd25685, 16'd23235, 16'd40016, 16'd17885, 16'd26676, 16'd1022, 16'd4643, 16'd54412, 16'd23506}; // indx = 307
    #10;
    addra = 32'd9856;
    dina = {96'd0, 16'd55918, 16'd35566, 16'd58525, 16'd11121, 16'd41300, 16'd4966, 16'd46113, 16'd9835, 16'd34233, 16'd31385}; // indx = 308
    #10;
    addra = 32'd9888;
    dina = {96'd0, 16'd14544, 16'd16337, 16'd48884, 16'd60558, 16'd43966, 16'd8806, 16'd15078, 16'd25016, 16'd43747, 16'd8929}; // indx = 309
    #10;
    addra = 32'd9920;
    dina = {96'd0, 16'd59127, 16'd12118, 16'd8260, 16'd7861, 16'd16036, 16'd41180, 16'd17669, 16'd41699, 16'd42055, 16'd32127}; // indx = 310
    #10;
    addra = 32'd9952;
    dina = {96'd0, 16'd46199, 16'd60150, 16'd42908, 16'd6790, 16'd63976, 16'd15397, 16'd63000, 16'd30614, 16'd32104, 16'd58509}; // indx = 311
    #10;
    addra = 32'd9984;
    dina = {96'd0, 16'd39807, 16'd33695, 16'd1803, 16'd29695, 16'd52472, 16'd1903, 16'd29562, 16'd13663, 16'd16988, 16'd27525}; // indx = 312
    #10;
    addra = 32'd10016;
    dina = {96'd0, 16'd13430, 16'd42980, 16'd24570, 16'd1101, 16'd50343, 16'd62632, 16'd21350, 16'd60235, 16'd41498, 16'd56233}; // indx = 313
    #10;
    addra = 32'd10048;
    dina = {96'd0, 16'd64703, 16'd13312, 16'd60917, 16'd34551, 16'd65227, 16'd61035, 16'd49045, 16'd41749, 16'd45873, 16'd4625}; // indx = 314
    #10;
    addra = 32'd10080;
    dina = {96'd0, 16'd23449, 16'd29164, 16'd46675, 16'd16748, 16'd41012, 16'd49508, 16'd6157, 16'd52150, 16'd13239, 16'd37668}; // indx = 315
    #10;
    addra = 32'd10112;
    dina = {96'd0, 16'd20346, 16'd59404, 16'd11543, 16'd64524, 16'd24186, 16'd22196, 16'd41154, 16'd61601, 16'd62047, 16'd34849}; // indx = 316
    #10;
    addra = 32'd10144;
    dina = {96'd0, 16'd26350, 16'd56603, 16'd60817, 16'd24779, 16'd4935, 16'd47956, 16'd27527, 16'd19296, 16'd33183, 16'd36908}; // indx = 317
    #10;
    addra = 32'd10176;
    dina = {96'd0, 16'd58104, 16'd25502, 16'd28200, 16'd21627, 16'd40713, 16'd18547, 16'd14314, 16'd50252, 16'd21246, 16'd33990}; // indx = 318
    #10;
    addra = 32'd10208;
    dina = {96'd0, 16'd62837, 16'd60597, 16'd52140, 16'd38849, 16'd24629, 16'd10952, 16'd36276, 16'd32244, 16'd506, 16'd36277}; // indx = 319
    #10;
    addra = 32'd10240;
    dina = {96'd0, 16'd18069, 16'd54510, 16'd32337, 16'd2048, 16'd46984, 16'd38380, 16'd27317, 16'd3119, 16'd43412, 16'd29984}; // indx = 320
    #10;
    addra = 32'd10272;
    dina = {96'd0, 16'd20177, 16'd60987, 16'd51070, 16'd48684, 16'd50713, 16'd44232, 16'd184, 16'd37001, 16'd31907, 16'd28198}; // indx = 321
    #10;
    addra = 32'd10304;
    dina = {96'd0, 16'd55339, 16'd36576, 16'd6641, 16'd440, 16'd56435, 16'd10041, 16'd34675, 16'd54439, 16'd3934, 16'd32531}; // indx = 322
    #10;
    addra = 32'd10336;
    dina = {96'd0, 16'd26919, 16'd11955, 16'd28298, 16'd26874, 16'd55906, 16'd55444, 16'd13554, 16'd64480, 16'd50820, 16'd34981}; // indx = 323
    #10;
    addra = 32'd10368;
    dina = {96'd0, 16'd19502, 16'd28270, 16'd52641, 16'd18932, 16'd53705, 16'd58166, 16'd10145, 16'd7328, 16'd43526, 16'd61139}; // indx = 324
    #10;
    addra = 32'd10400;
    dina = {96'd0, 16'd23925, 16'd32456, 16'd27329, 16'd1708, 16'd38388, 16'd59063, 16'd26075, 16'd44429, 16'd9859, 16'd52436}; // indx = 325
    #10;
    addra = 32'd10432;
    dina = {96'd0, 16'd12081, 16'd6325, 16'd59658, 16'd20997, 16'd49987, 16'd25302, 16'd29359, 16'd48801, 16'd20701, 16'd52168}; // indx = 326
    #10;
    addra = 32'd10464;
    dina = {96'd0, 16'd36823, 16'd4348, 16'd11378, 16'd1051, 16'd56106, 16'd28332, 16'd42059, 16'd60552, 16'd11900, 16'd102}; // indx = 327
    #10;
    addra = 32'd10496;
    dina = {96'd0, 16'd49161, 16'd47190, 16'd35064, 16'd11193, 16'd5042, 16'd59684, 16'd51673, 16'd42810, 16'd38849, 16'd46043}; // indx = 328
    #10;
    addra = 32'd10528;
    dina = {96'd0, 16'd8101, 16'd20806, 16'd14212, 16'd18030, 16'd43610, 16'd41636, 16'd59380, 16'd31752, 16'd61969, 16'd9117}; // indx = 329
    #10;
    addra = 32'd10560;
    dina = {96'd0, 16'd14183, 16'd51976, 16'd60622, 16'd26786, 16'd59822, 16'd50787, 16'd42689, 16'd16801, 16'd18826, 16'd223}; // indx = 330
    #10;
    addra = 32'd10592;
    dina = {96'd0, 16'd43277, 16'd44083, 16'd62354, 16'd56647, 16'd59408, 16'd3756, 16'd5579, 16'd12486, 16'd46327, 16'd61995}; // indx = 331
    #10;
    addra = 32'd10624;
    dina = {96'd0, 16'd47749, 16'd45770, 16'd32295, 16'd45936, 16'd49272, 16'd21432, 16'd10566, 16'd54822, 16'd37197, 16'd32413}; // indx = 332
    #10;
    addra = 32'd10656;
    dina = {96'd0, 16'd25224, 16'd45300, 16'd39564, 16'd36853, 16'd8990, 16'd64589, 16'd43956, 16'd31977, 16'd13474, 16'd39274}; // indx = 333
    #10;
    addra = 32'd10688;
    dina = {96'd0, 16'd29043, 16'd43430, 16'd60396, 16'd51705, 16'd29012, 16'd62427, 16'd711, 16'd6347, 16'd11643, 16'd52834}; // indx = 334
    #10;
    addra = 32'd10720;
    dina = {96'd0, 16'd1468, 16'd43335, 16'd57388, 16'd11382, 16'd31105, 16'd25548, 16'd33045, 16'd43780, 16'd6575, 16'd42091}; // indx = 335
    #10;
    addra = 32'd10752;
    dina = {96'd0, 16'd47168, 16'd61827, 16'd64736, 16'd27047, 16'd58766, 16'd6684, 16'd25262, 16'd19458, 16'd55383, 16'd50826}; // indx = 336
    #10;
    addra = 32'd10784;
    dina = {96'd0, 16'd62906, 16'd5073, 16'd52986, 16'd15746, 16'd21811, 16'd44126, 16'd59743, 16'd65150, 16'd58746, 16'd56067}; // indx = 337
    #10;
    addra = 32'd10816;
    dina = {96'd0, 16'd30790, 16'd4889, 16'd25869, 16'd17011, 16'd8962, 16'd36275, 16'd52043, 16'd49147, 16'd62581, 16'd27689}; // indx = 338
    #10;
    addra = 32'd10848;
    dina = {96'd0, 16'd13342, 16'd45571, 16'd40278, 16'd60390, 16'd44549, 16'd56287, 16'd55715, 16'd18419, 16'd43500, 16'd6359}; // indx = 339
    #10;
    addra = 32'd10880;
    dina = {96'd0, 16'd42152, 16'd23257, 16'd57534, 16'd59108, 16'd27301, 16'd6576, 16'd19142, 16'd21946, 16'd35154, 16'd26443}; // indx = 340
    #10;
    addra = 32'd10912;
    dina = {96'd0, 16'd29121, 16'd44205, 16'd2351, 16'd6352, 16'd48954, 16'd40653, 16'd20480, 16'd23584, 16'd40130, 16'd13733}; // indx = 341
    #10;
    addra = 32'd10944;
    dina = {96'd0, 16'd7811, 16'd28781, 16'd52423, 16'd21605, 16'd26879, 16'd11471, 16'd10122, 16'd11419, 16'd41356, 16'd29532}; // indx = 342
    #10;
    addra = 32'd10976;
    dina = {96'd0, 16'd53906, 16'd12154, 16'd15485, 16'd19159, 16'd1120, 16'd10911, 16'd24912, 16'd10542, 16'd8753, 16'd1600}; // indx = 343
    #10;
    addra = 32'd11008;
    dina = {96'd0, 16'd46340, 16'd43258, 16'd17729, 16'd63806, 16'd39303, 16'd42534, 16'd21523, 16'd9137, 16'd37542, 16'd64426}; // indx = 344
    #10;
    addra = 32'd11040;
    dina = {96'd0, 16'd42767, 16'd56006, 16'd22164, 16'd9847, 16'd51610, 16'd19507, 16'd63185, 16'd55302, 16'd14914, 16'd58142}; // indx = 345
    #10;
    addra = 32'd11072;
    dina = {96'd0, 16'd59014, 16'd8628, 16'd7513, 16'd1793, 16'd51019, 16'd47462, 16'd23781, 16'd39891, 16'd8876, 16'd50307}; // indx = 346
    #10;
    addra = 32'd11104;
    dina = {96'd0, 16'd57225, 16'd29265, 16'd6852, 16'd28455, 16'd35656, 16'd11001, 16'd58897, 16'd23118, 16'd49571, 16'd59403}; // indx = 347
    #10;
    addra = 32'd11136;
    dina = {96'd0, 16'd1144, 16'd64049, 16'd39984, 16'd47428, 16'd37247, 16'd4426, 16'd47252, 16'd7830, 16'd36839, 16'd52615}; // indx = 348
    #10;
    addra = 32'd11168;
    dina = {96'd0, 16'd40868, 16'd49028, 16'd24354, 16'd1862, 16'd31096, 16'd62920, 16'd18911, 16'd21314, 16'd18071, 16'd56498}; // indx = 349
    #10;
    addra = 32'd11200;
    dina = {96'd0, 16'd55792, 16'd7003, 16'd41552, 16'd52206, 16'd2892, 16'd18914, 16'd46772, 16'd54301, 16'd65288, 16'd13183}; // indx = 350
    #10;
    addra = 32'd11232;
    dina = {96'd0, 16'd2095, 16'd5472, 16'd27257, 16'd6797, 16'd37615, 16'd51104, 16'd37629, 16'd32447, 16'd53968, 16'd26797}; // indx = 351
    #10;
    addra = 32'd11264;
    dina = {96'd0, 16'd11203, 16'd21556, 16'd9965, 16'd65228, 16'd4184, 16'd54655, 16'd61956, 16'd21766, 16'd29017, 16'd13904}; // indx = 352
    #10;
    addra = 32'd11296;
    dina = {96'd0, 16'd60958, 16'd31504, 16'd5041, 16'd8165, 16'd18805, 16'd13377, 16'd57692, 16'd34246, 16'd330, 16'd43916}; // indx = 353
    #10;
    addra = 32'd11328;
    dina = {96'd0, 16'd3501, 16'd33695, 16'd47073, 16'd51096, 16'd1652, 16'd40849, 16'd47691, 16'd17799, 16'd31301, 16'd11138}; // indx = 354
    #10;
    addra = 32'd11360;
    dina = {96'd0, 16'd48884, 16'd37432, 16'd55467, 16'd55231, 16'd49234, 16'd63393, 16'd52895, 16'd51383, 16'd4710, 16'd8209}; // indx = 355
    #10;
    addra = 32'd11392;
    dina = {96'd0, 16'd62915, 16'd51046, 16'd38401, 16'd22502, 16'd11231, 16'd4994, 16'd10212, 16'd42234, 16'd7000, 16'd46790}; // indx = 356
    #10;
    addra = 32'd11424;
    dina = {96'd0, 16'd22489, 16'd26916, 16'd56614, 16'd4161, 16'd57665, 16'd18067, 16'd24802, 16'd39474, 16'd7406, 16'd28153}; // indx = 357
    #10;
    addra = 32'd11456;
    dina = {96'd0, 16'd50519, 16'd9455, 16'd5640, 16'd6865, 16'd38409, 16'd7368, 16'd64725, 16'd8673, 16'd26685, 16'd1520}; // indx = 358
    #10;
    addra = 32'd11488;
    dina = {96'd0, 16'd28854, 16'd45439, 16'd18375, 16'd16190, 16'd5329, 16'd4464, 16'd54873, 16'd45983, 16'd13162, 16'd15358}; // indx = 359
    #10;
    addra = 32'd11520;
    dina = {96'd0, 16'd20058, 16'd28576, 16'd16390, 16'd17049, 16'd64551, 16'd35386, 16'd20846, 16'd16051, 16'd4117, 16'd8305}; // indx = 360
    #10;
    addra = 32'd11552;
    dina = {96'd0, 16'd19466, 16'd40662, 16'd10018, 16'd20452, 16'd61003, 16'd37284, 16'd62482, 16'd2835, 16'd8002, 16'd40735}; // indx = 361
    #10;
    addra = 32'd11584;
    dina = {96'd0, 16'd48117, 16'd14572, 16'd27729, 16'd64714, 16'd47739, 16'd325, 16'd38880, 16'd9765, 16'd5957, 16'd58944}; // indx = 362
    #10;
    addra = 32'd11616;
    dina = {96'd0, 16'd22170, 16'd30580, 16'd59636, 16'd60797, 16'd20094, 16'd58962, 16'd39904, 16'd29380, 16'd29453, 16'd64217}; // indx = 363
    #10;
    addra = 32'd11648;
    dina = {96'd0, 16'd16214, 16'd31784, 16'd52624, 16'd35405, 16'd19415, 16'd61804, 16'd39803, 16'd5898, 16'd61322, 16'd13064}; // indx = 364
    #10;
    addra = 32'd11680;
    dina = {96'd0, 16'd49682, 16'd58098, 16'd51824, 16'd3890, 16'd10902, 16'd20810, 16'd51982, 16'd32421, 16'd28160, 16'd40261}; // indx = 365
    #10;
    addra = 32'd11712;
    dina = {96'd0, 16'd23521, 16'd40660, 16'd10488, 16'd12408, 16'd28042, 16'd20128, 16'd28258, 16'd35844, 16'd9388, 16'd25738}; // indx = 366
    #10;
    addra = 32'd11744;
    dina = {96'd0, 16'd11605, 16'd24457, 16'd44999, 16'd44254, 16'd8104, 16'd43696, 16'd35122, 16'd20950, 16'd40508, 16'd64454}; // indx = 367
    #10;
    addra = 32'd11776;
    dina = {96'd0, 16'd39839, 16'd23268, 16'd59678, 16'd13038, 16'd31170, 16'd56194, 16'd577, 16'd20848, 16'd14560, 16'd28301}; // indx = 368
    #10;
    addra = 32'd11808;
    dina = {96'd0, 16'd44757, 16'd31642, 16'd42188, 16'd63044, 16'd51635, 16'd12970, 16'd11748, 16'd49626, 16'd44154, 16'd17191}; // indx = 369
    #10;
    addra = 32'd11840;
    dina = {96'd0, 16'd13030, 16'd56474, 16'd6090, 16'd7991, 16'd20619, 16'd2658, 16'd56117, 16'd19148, 16'd60045, 16'd23265}; // indx = 370
    #10;
    addra = 32'd11872;
    dina = {96'd0, 16'd37718, 16'd46888, 16'd30110, 16'd28677, 16'd14656, 16'd45047, 16'd4833, 16'd58437, 16'd65182, 16'd1689}; // indx = 371
    #10;
    addra = 32'd11904;
    dina = {96'd0, 16'd64529, 16'd43301, 16'd32274, 16'd27475, 16'd63202, 16'd3683, 16'd48731, 16'd27580, 16'd27900, 16'd22468}; // indx = 372
    #10;
    addra = 32'd11936;
    dina = {96'd0, 16'd48998, 16'd22331, 16'd43734, 16'd20610, 16'd15012, 16'd5220, 16'd54250, 16'd12143, 16'd38971, 16'd42800}; // indx = 373
    #10;
    addra = 32'd11968;
    dina = {96'd0, 16'd26381, 16'd64829, 16'd11375, 16'd59552, 16'd16245, 16'd25019, 16'd49630, 16'd51565, 16'd22279, 16'd5698}; // indx = 374
    #10;
    addra = 32'd12000;
    dina = {96'd0, 16'd48712, 16'd27010, 16'd45222, 16'd39105, 16'd59560, 16'd28045, 16'd15693, 16'd41148, 16'd36045, 16'd60177}; // indx = 375
    #10;
    addra = 32'd12032;
    dina = {96'd0, 16'd21337, 16'd23555, 16'd45820, 16'd24858, 16'd13685, 16'd11258, 16'd4494, 16'd21471, 16'd63889, 16'd25839}; // indx = 376
    #10;
    addra = 32'd12064;
    dina = {96'd0, 16'd8990, 16'd46175, 16'd31784, 16'd575, 16'd63674, 16'd26185, 16'd6258, 16'd21010, 16'd14989, 16'd55757}; // indx = 377
    #10;
    addra = 32'd12096;
    dina = {96'd0, 16'd46703, 16'd52373, 16'd36968, 16'd11295, 16'd34975, 16'd56275, 16'd59947, 16'd54015, 16'd63037, 16'd31820}; // indx = 378
    #10;
    addra = 32'd12128;
    dina = {96'd0, 16'd50819, 16'd30327, 16'd40810, 16'd12535, 16'd30134, 16'd15406, 16'd55406, 16'd32828, 16'd6208, 16'd59248}; // indx = 379
    #10;
    addra = 32'd12160;
    dina = {96'd0, 16'd24811, 16'd46612, 16'd6843, 16'd28262, 16'd47621, 16'd18155, 16'd38650, 16'd49399, 16'd64957, 16'd63700}; // indx = 380
    #10;
    addra = 32'd12192;
    dina = {96'd0, 16'd21866, 16'd37006, 16'd26107, 16'd25168, 16'd54326, 16'd7586, 16'd41029, 16'd50602, 16'd62245, 16'd18905}; // indx = 381
    #10;
    addra = 32'd12224;
    dina = {96'd0, 16'd57757, 16'd17103, 16'd34587, 16'd22555, 16'd15491, 16'd24664, 16'd28319, 16'd41638, 16'd55552, 16'd11311}; // indx = 382
    #10;
    addra = 32'd12256;
    dina = {96'd0, 16'd37349, 16'd55639, 16'd31642, 16'd41091, 16'd35596, 16'd47842, 16'd53089, 16'd2975, 16'd10918, 16'd52888}; // indx = 383
    #10;
    addra = 32'd12288;
    dina = {96'd0, 16'd36845, 16'd31805, 16'd34940, 16'd11192, 16'd49728, 16'd2129, 16'd55632, 16'd4732, 16'd23134, 16'd5}; // indx = 384
    #10;
    addra = 32'd12320;
    dina = {96'd0, 16'd52251, 16'd8328, 16'd24606, 16'd56863, 16'd16348, 16'd32513, 16'd49077, 16'd46483, 16'd6142, 16'd6273}; // indx = 385
    #10;
    addra = 32'd12352;
    dina = {96'd0, 16'd4571, 16'd54948, 16'd65345, 16'd13897, 16'd24842, 16'd44810, 16'd41050, 16'd24440, 16'd16469, 16'd28169}; // indx = 386
    #10;
    addra = 32'd12384;
    dina = {96'd0, 16'd31655, 16'd52754, 16'd45715, 16'd52843, 16'd19219, 16'd27716, 16'd17492, 16'd2063, 16'd2237, 16'd21458}; // indx = 387
    #10;
    addra = 32'd12416;
    dina = {96'd0, 16'd23780, 16'd43604, 16'd31574, 16'd26580, 16'd27897, 16'd13681, 16'd59125, 16'd20036, 16'd20486, 16'd20320}; // indx = 388
    #10;
    addra = 32'd12448;
    dina = {96'd0, 16'd48848, 16'd59099, 16'd4328, 16'd25619, 16'd14969, 16'd11153, 16'd44623, 16'd35440, 16'd39462, 16'd41479}; // indx = 389
    #10;
    addra = 32'd12480;
    dina = {96'd0, 16'd1703, 16'd27376, 16'd6887, 16'd22192, 16'd35072, 16'd23311, 16'd14200, 16'd42196, 16'd4677, 16'd22347}; // indx = 390
    #10;
    addra = 32'd12512;
    dina = {96'd0, 16'd5357, 16'd15946, 16'd62355, 16'd23024, 16'd3867, 16'd58142, 16'd46054, 16'd6522, 16'd26251, 16'd36606}; // indx = 391
    #10;
    addra = 32'd12544;
    dina = {96'd0, 16'd13060, 16'd50156, 16'd13110, 16'd19039, 16'd26793, 16'd10833, 16'd60153, 16'd27833, 16'd24497, 16'd2452}; // indx = 392
    #10;
    addra = 32'd12576;
    dina = {96'd0, 16'd13499, 16'd48574, 16'd31141, 16'd29530, 16'd55782, 16'd10019, 16'd11164, 16'd41276, 16'd58165, 16'd63422}; // indx = 393
    #10;
    addra = 32'd12608;
    dina = {96'd0, 16'd49147, 16'd33727, 16'd28757, 16'd18597, 16'd51519, 16'd23657, 16'd22649, 16'd52803, 16'd28580, 16'd15932}; // indx = 394
    #10;
    addra = 32'd12640;
    dina = {96'd0, 16'd2896, 16'd49810, 16'd31649, 16'd13074, 16'd32868, 16'd9275, 16'd45411, 16'd36423, 16'd33905, 16'd22191}; // indx = 395
    #10;
    addra = 32'd12672;
    dina = {96'd0, 16'd47772, 16'd25826, 16'd32633, 16'd36202, 16'd34123, 16'd19814, 16'd22628, 16'd34967, 16'd39174, 16'd18931}; // indx = 396
    #10;
    addra = 32'd12704;
    dina = {96'd0, 16'd20778, 16'd23734, 16'd62113, 16'd6084, 16'd34864, 16'd40996, 16'd30261, 16'd38317, 16'd4459, 16'd65207}; // indx = 397
    #10;
    addra = 32'd12736;
    dina = {96'd0, 16'd21380, 16'd37791, 16'd7304, 16'd5227, 16'd43518, 16'd803, 16'd29557, 16'd42536, 16'd28792, 16'd28000}; // indx = 398
    #10;
    addra = 32'd12768;
    dina = {96'd0, 16'd17638, 16'd63794, 16'd31227, 16'd33177, 16'd6042, 16'd18907, 16'd36120, 16'd58311, 16'd38302, 16'd6628}; // indx = 399
    #10;
    addra = 32'd12800;
    dina = {96'd0, 16'd14375, 16'd35131, 16'd28550, 16'd24283, 16'd24601, 16'd48111, 16'd42628, 16'd16642, 16'd16368, 16'd16983}; // indx = 400
    #10;
    addra = 32'd12832;
    dina = {96'd0, 16'd54649, 16'd41885, 16'd1638, 16'd50720, 16'd59790, 16'd8746, 16'd65452, 16'd24710, 16'd60033, 16'd32767}; // indx = 401
    #10;
    addra = 32'd12864;
    dina = {96'd0, 16'd16354, 16'd1087, 16'd58991, 16'd65192, 16'd20573, 16'd18285, 16'd36408, 16'd18931, 16'd12293, 16'd49026}; // indx = 402
    #10;
    addra = 32'd12896;
    dina = {96'd0, 16'd6270, 16'd39794, 16'd708, 16'd63457, 16'd4110, 16'd39688, 16'd6344, 16'd2402, 16'd62174, 16'd7190}; // indx = 403
    #10;
    addra = 32'd12928;
    dina = {96'd0, 16'd25817, 16'd46701, 16'd61217, 16'd55419, 16'd56874, 16'd44661, 16'd26519, 16'd18298, 16'd33424, 16'd11887}; // indx = 404
    #10;
    addra = 32'd12960;
    dina = {96'd0, 16'd25452, 16'd38088, 16'd49180, 16'd1977, 16'd56172, 16'd19690, 16'd36770, 16'd37813, 16'd21575, 16'd47945}; // indx = 405
    #10;
    addra = 32'd12992;
    dina = {96'd0, 16'd2468, 16'd54023, 16'd37013, 16'd21705, 16'd36548, 16'd57999, 16'd34737, 16'd7859, 16'd11055, 16'd14313}; // indx = 406
    #10;
    addra = 32'd13024;
    dina = {96'd0, 16'd10373, 16'd38211, 16'd2061, 16'd59158, 16'd43239, 16'd43628, 16'd59646, 16'd64624, 16'd22241, 16'd18270}; // indx = 407
    #10;
    addra = 32'd13056;
    dina = {96'd0, 16'd15836, 16'd64084, 16'd57439, 16'd47020, 16'd6132, 16'd29059, 16'd47192, 16'd32, 16'd18454, 16'd55796}; // indx = 408
    #10;
    addra = 32'd13088;
    dina = {96'd0, 16'd63753, 16'd42004, 16'd56888, 16'd21757, 16'd9312, 16'd41897, 16'd13900, 16'd61971, 16'd30554, 16'd679}; // indx = 409
    #10;
    addra = 32'd13120;
    dina = {96'd0, 16'd65064, 16'd45542, 16'd21452, 16'd9494, 16'd7724, 16'd62633, 16'd37456, 16'd2397, 16'd60294, 16'd24232}; // indx = 410
    #10;
    addra = 32'd13152;
    dina = {96'd0, 16'd30117, 16'd3197, 16'd10606, 16'd33392, 16'd3500, 16'd41381, 16'd50580, 16'd1132, 16'd10844, 16'd36029}; // indx = 411
    #10;
    addra = 32'd13184;
    dina = {96'd0, 16'd866, 16'd42933, 16'd56591, 16'd56069, 16'd45839, 16'd51500, 16'd50861, 16'd33791, 16'd39196, 16'd46985}; // indx = 412
    #10;
    addra = 32'd13216;
    dina = {96'd0, 16'd41164, 16'd17729, 16'd20555, 16'd10057, 16'd48993, 16'd60251, 16'd50976, 16'd15871, 16'd52953, 16'd34330}; // indx = 413
    #10;
    addra = 32'd13248;
    dina = {96'd0, 16'd62809, 16'd2903, 16'd4647, 16'd35650, 16'd21493, 16'd60509, 16'd32808, 16'd6900, 16'd23126, 16'd60595}; // indx = 414
    #10;
    addra = 32'd13280;
    dina = {96'd0, 16'd21046, 16'd56177, 16'd43980, 16'd19987, 16'd30764, 16'd23016, 16'd27270, 16'd38556, 16'd9549, 16'd55555}; // indx = 415
    #10;
    addra = 32'd13312;
    dina = {96'd0, 16'd62938, 16'd27922, 16'd55465, 16'd26761, 16'd51765, 16'd19419, 16'd61087, 16'd12067, 16'd26345, 16'd5819}; // indx = 416
    #10;
    addra = 32'd13344;
    dina = {96'd0, 16'd51908, 16'd46570, 16'd18667, 16'd23406, 16'd12064, 16'd45353, 16'd10983, 16'd18282, 16'd10125, 16'd39462}; // indx = 417
    #10;
    addra = 32'd13376;
    dina = {96'd0, 16'd45238, 16'd45847, 16'd39339, 16'd42413, 16'd56300, 16'd60588, 16'd41409, 16'd8208, 16'd24827, 16'd44839}; // indx = 418
    #10;
    addra = 32'd13408;
    dina = {96'd0, 16'd52936, 16'd63895, 16'd60366, 16'd9812, 16'd18453, 16'd22087, 16'd43903, 16'd53358, 16'd29855, 16'd37234}; // indx = 419
    #10;
    addra = 32'd13440;
    dina = {96'd0, 16'd63877, 16'd51746, 16'd18977, 16'd56475, 16'd164, 16'd37457, 16'd32812, 16'd11086, 16'd43143, 16'd45786}; // indx = 420
    #10;
    addra = 32'd13472;
    dina = {96'd0, 16'd22498, 16'd38857, 16'd56147, 16'd41873, 16'd16540, 16'd23390, 16'd17148, 16'd60474, 16'd57054, 16'd52029}; // indx = 421
    #10;
    addra = 32'd13504;
    dina = {96'd0, 16'd9009, 16'd36876, 16'd64847, 16'd16684, 16'd25023, 16'd55508, 16'd11661, 16'd65287, 16'd8480, 16'd39458}; // indx = 422
    #10;
    addra = 32'd13536;
    dina = {96'd0, 16'd59289, 16'd7143, 16'd43582, 16'd49707, 16'd35096, 16'd60808, 16'd12215, 16'd57049, 16'd54645, 16'd27719}; // indx = 423
    #10;
    addra = 32'd13568;
    dina = {96'd0, 16'd47653, 16'd10846, 16'd37922, 16'd40607, 16'd25736, 16'd45858, 16'd22506, 16'd44967, 16'd14374, 16'd18697}; // indx = 424
    #10;
    addra = 32'd13600;
    dina = {96'd0, 16'd46094, 16'd31349, 16'd35259, 16'd60039, 16'd54072, 16'd34239, 16'd3509, 16'd55131, 16'd62827, 16'd44681}; // indx = 425
    #10;
    addra = 32'd13632;
    dina = {96'd0, 16'd37804, 16'd59881, 16'd38018, 16'd4473, 16'd49363, 16'd10969, 16'd32573, 16'd45028, 16'd21650, 16'd2576}; // indx = 426
    #10;
    addra = 32'd13664;
    dina = {96'd0, 16'd27068, 16'd35045, 16'd6808, 16'd15842, 16'd37224, 16'd20283, 16'd42448, 16'd12862, 16'd48712, 16'd50765}; // indx = 427
    #10;
    addra = 32'd13696;
    dina = {96'd0, 16'd4148, 16'd6280, 16'd4758, 16'd18950, 16'd37032, 16'd32617, 16'd15461, 16'd36496, 16'd37561, 16'd7049}; // indx = 428
    #10;
    addra = 32'd13728;
    dina = {96'd0, 16'd14545, 16'd48897, 16'd50149, 16'd49609, 16'd2769, 16'd15652, 16'd32871, 16'd9630, 16'd36426, 16'd42904}; // indx = 429
    #10;
    addra = 32'd13760;
    dina = {96'd0, 16'd58560, 16'd51848, 16'd4683, 16'd62885, 16'd14775, 16'd24450, 16'd757, 16'd45630, 16'd27228, 16'd11609}; // indx = 430
    #10;
    addra = 32'd13792;
    dina = {96'd0, 16'd65097, 16'd14204, 16'd33838, 16'd43166, 16'd23786, 16'd50569, 16'd11199, 16'd6150, 16'd41396, 16'd11419}; // indx = 431
    #10;
    addra = 32'd13824;
    dina = {96'd0, 16'd54376, 16'd63141, 16'd26662, 16'd18780, 16'd8331, 16'd1529, 16'd63762, 16'd4115, 16'd17312, 16'd55561}; // indx = 432
    #10;
    addra = 32'd13856;
    dina = {96'd0, 16'd55089, 16'd63574, 16'd21242, 16'd33304, 16'd3486, 16'd36214, 16'd43421, 16'd58390, 16'd62941, 16'd24163}; // indx = 433
    #10;
    addra = 32'd13888;
    dina = {96'd0, 16'd41786, 16'd52648, 16'd31308, 16'd33071, 16'd12934, 16'd57413, 16'd64515, 16'd5929, 16'd56621, 16'd33977}; // indx = 434
    #10;
    addra = 32'd13920;
    dina = {96'd0, 16'd422, 16'd33959, 16'd16683, 16'd26471, 16'd63229, 16'd28182, 16'd6163, 16'd1653, 16'd61929, 16'd30683}; // indx = 435
    #10;
    addra = 32'd13952;
    dina = {96'd0, 16'd42812, 16'd50117, 16'd63841, 16'd64498, 16'd15287, 16'd64410, 16'd47587, 16'd19665, 16'd64048, 16'd49127}; // indx = 436
    #10;
    addra = 32'd13984;
    dina = {96'd0, 16'd35467, 16'd28541, 16'd6517, 16'd48536, 16'd61047, 16'd881, 16'd41879, 16'd43838, 16'd7705, 16'd47132}; // indx = 437
    #10;
    addra = 32'd14016;
    dina = {96'd0, 16'd29651, 16'd9464, 16'd55756, 16'd3537, 16'd28843, 16'd45596, 16'd46416, 16'd45600, 16'd4726, 16'd56804}; // indx = 438
    #10;
    addra = 32'd14048;
    dina = {96'd0, 16'd14389, 16'd7562, 16'd6681, 16'd22881, 16'd42126, 16'd59151, 16'd7709, 16'd57099, 16'd48816, 16'd3385}; // indx = 439
    #10;
    addra = 32'd14080;
    dina = {96'd0, 16'd11903, 16'd58275, 16'd34974, 16'd2746, 16'd4019, 16'd46413, 16'd23704, 16'd40064, 16'd11068, 16'd52702}; // indx = 440
    #10;
    addra = 32'd14112;
    dina = {96'd0, 16'd23852, 16'd35415, 16'd42440, 16'd38387, 16'd2082, 16'd56058, 16'd54130, 16'd17105, 16'd55463, 16'd42332}; // indx = 441
    #10;
    addra = 32'd14144;
    dina = {96'd0, 16'd54898, 16'd46272, 16'd37978, 16'd31699, 16'd35874, 16'd16232, 16'd37441, 16'd56125, 16'd50128, 16'd58422}; // indx = 442
    #10;
    addra = 32'd14176;
    dina = {96'd0, 16'd32465, 16'd20422, 16'd37048, 16'd22485, 16'd50674, 16'd35971, 16'd46735, 16'd4048, 16'd64513, 16'd65401}; // indx = 443
    #10;
    addra = 32'd14208;
    dina = {96'd0, 16'd22617, 16'd29912, 16'd48213, 16'd62432, 16'd13170, 16'd17034, 16'd50975, 16'd34462, 16'd19491, 16'd59646}; // indx = 444
    #10;
    addra = 32'd14240;
    dina = {96'd0, 16'd63962, 16'd23255, 16'd36218, 16'd1751, 16'd33326, 16'd47449, 16'd27013, 16'd24923, 16'd13624, 16'd29425}; // indx = 445
    #10;
    addra = 32'd14272;
    dina = {96'd0, 16'd27736, 16'd53551, 16'd12789, 16'd22046, 16'd52121, 16'd50776, 16'd42143, 16'd30906, 16'd53014, 16'd17420}; // indx = 446
    #10;
    addra = 32'd14304;
    dina = {96'd0, 16'd12677, 16'd50696, 16'd28528, 16'd11611, 16'd40352, 16'd27396, 16'd64160, 16'd30487, 16'd24043, 16'd21599}; // indx = 447
    #10;
    addra = 32'd14336;
    dina = {96'd0, 16'd54569, 16'd16243, 16'd9793, 16'd49783, 16'd36199, 16'd25721, 16'd37135, 16'd26150, 16'd49092, 16'd20905}; // indx = 448
    #10;
    addra = 32'd14368;
    dina = {96'd0, 16'd64254, 16'd25984, 16'd11070, 16'd16793, 16'd63384, 16'd29458, 16'd34297, 16'd19638, 16'd39615, 16'd35596}; // indx = 449
    #10;
    addra = 32'd14400;
    dina = {96'd0, 16'd20955, 16'd44350, 16'd39456, 16'd39014, 16'd12793, 16'd7744, 16'd7868, 16'd57990, 16'd58751, 16'd18069}; // indx = 450
    #10;
    addra = 32'd14432;
    dina = {96'd0, 16'd56789, 16'd35866, 16'd6025, 16'd26254, 16'd35482, 16'd57250, 16'd33003, 16'd37074, 16'd25537, 16'd44275}; // indx = 451
    #10;
    addra = 32'd14464;
    dina = {96'd0, 16'd60579, 16'd46061, 16'd18673, 16'd61127, 16'd6330, 16'd57712, 16'd7383, 16'd57193, 16'd61028, 16'd54773}; // indx = 452
    #10;
    addra = 32'd14496;
    dina = {96'd0, 16'd47921, 16'd51113, 16'd7797, 16'd1464, 16'd1285, 16'd56737, 16'd62472, 16'd63398, 16'd52234, 16'd50650}; // indx = 453
    #10;
    addra = 32'd14528;
    dina = {96'd0, 16'd8024, 16'd15384, 16'd9247, 16'd38782, 16'd38711, 16'd60152, 16'd53779, 16'd526, 16'd52936, 16'd28407}; // indx = 454
    #10;
    addra = 32'd14560;
    dina = {96'd0, 16'd42720, 16'd24209, 16'd45317, 16'd58116, 16'd58942, 16'd43518, 16'd27719, 16'd43416, 16'd13831, 16'd51832}; // indx = 455
    #10;
    addra = 32'd14592;
    dina = {96'd0, 16'd58616, 16'd19406, 16'd37535, 16'd4188, 16'd64209, 16'd18354, 16'd41432, 16'd63234, 16'd2606, 16'd24553}; // indx = 456
    #10;
    addra = 32'd14624;
    dina = {96'd0, 16'd31982, 16'd51542, 16'd33068, 16'd46737, 16'd7904, 16'd37482, 16'd17830, 16'd50743, 16'd54120, 16'd27681}; // indx = 457
    #10;
    addra = 32'd14656;
    dina = {96'd0, 16'd57197, 16'd42649, 16'd63389, 16'd39871, 16'd54874, 16'd46753, 16'd29144, 16'd54229, 16'd36955, 16'd19522}; // indx = 458
    #10;
    addra = 32'd14688;
    dina = {96'd0, 16'd23660, 16'd4111, 16'd58660, 16'd16649, 16'd16051, 16'd60097, 16'd42073, 16'd8490, 16'd25624, 16'd37947}; // indx = 459
    #10;
    addra = 32'd14720;
    dina = {96'd0, 16'd17766, 16'd62554, 16'd14835, 16'd48866, 16'd56684, 16'd62789, 16'd37618, 16'd1891, 16'd59948, 16'd41563}; // indx = 460
    #10;
    addra = 32'd14752;
    dina = {96'd0, 16'd37104, 16'd52653, 16'd29609, 16'd39397, 16'd65179, 16'd25032, 16'd21078, 16'd33929, 16'd43117, 16'd19439}; // indx = 461
    #10;
    addra = 32'd14784;
    dina = {96'd0, 16'd39821, 16'd828, 16'd13839, 16'd47782, 16'd13014, 16'd1486, 16'd17195, 16'd9568, 16'd23233, 16'd19547}; // indx = 462
    #10;
    addra = 32'd14816;
    dina = {96'd0, 16'd49200, 16'd65054, 16'd522, 16'd33997, 16'd44962, 16'd24217, 16'd54386, 16'd59732, 16'd49478, 16'd15063}; // indx = 463
    #10;
    addra = 32'd14848;
    dina = {96'd0, 16'd22942, 16'd29304, 16'd27670, 16'd24524, 16'd53594, 16'd956, 16'd58038, 16'd52534, 16'd32030, 16'd51142}; // indx = 464
    #10;
    addra = 32'd14880;
    dina = {96'd0, 16'd36260, 16'd61261, 16'd17827, 16'd11084, 16'd47015, 16'd65064, 16'd55566, 16'd21185, 16'd24517, 16'd37605}; // indx = 465
    #10;
    addra = 32'd14912;
    dina = {96'd0, 16'd64762, 16'd18169, 16'd63338, 16'd65003, 16'd17658, 16'd51778, 16'd44355, 16'd42499, 16'd45147, 16'd4023}; // indx = 466
    #10;
    addra = 32'd14944;
    dina = {96'd0, 16'd64297, 16'd56590, 16'd35241, 16'd10375, 16'd53340, 16'd5811, 16'd3736, 16'd49911, 16'd19165, 16'd56990}; // indx = 467
    #10;
    addra = 32'd14976;
    dina = {96'd0, 16'd46043, 16'd27100, 16'd51188, 16'd25690, 16'd25146, 16'd42457, 16'd50047, 16'd32913, 16'd30144, 16'd62402}; // indx = 468
    #10;
    addra = 32'd15008;
    dina = {96'd0, 16'd21694, 16'd65258, 16'd27569, 16'd16323, 16'd28827, 16'd56112, 16'd3773, 16'd56947, 16'd13021, 16'd24153}; // indx = 469
    #10;
    addra = 32'd15040;
    dina = {96'd0, 16'd20482, 16'd35198, 16'd52002, 16'd51391, 16'd60300, 16'd53656, 16'd36123, 16'd1556, 16'd28002, 16'd47589}; // indx = 470
    #10;
    addra = 32'd15072;
    dina = {96'd0, 16'd38441, 16'd38765, 16'd54372, 16'd43583, 16'd1644, 16'd52336, 16'd35244, 16'd52360, 16'd8747, 16'd47989}; // indx = 471
    #10;
    addra = 32'd15104;
    dina = {96'd0, 16'd34395, 16'd56751, 16'd12779, 16'd59698, 16'd9509, 16'd3307, 16'd28456, 16'd48407, 16'd33252, 16'd2105}; // indx = 472
    #10;
    addra = 32'd15136;
    dina = {96'd0, 16'd26899, 16'd11175, 16'd33565, 16'd26836, 16'd61466, 16'd26037, 16'd1101, 16'd39389, 16'd28275, 16'd23152}; // indx = 473
    #10;
    addra = 32'd15168;
    dina = {96'd0, 16'd59435, 16'd2357, 16'd39732, 16'd31347, 16'd39384, 16'd51659, 16'd61131, 16'd53056, 16'd46672, 16'd53595}; // indx = 474
    #10;
    addra = 32'd15200;
    dina = {96'd0, 16'd40815, 16'd18293, 16'd1444, 16'd49809, 16'd37998, 16'd63822, 16'd29365, 16'd35999, 16'd3708, 16'd47070}; // indx = 475
    #10;
    addra = 32'd15232;
    dina = {96'd0, 16'd51259, 16'd8233, 16'd61119, 16'd28125, 16'd413, 16'd48471, 16'd8069, 16'd60248, 16'd57236, 16'd11655}; // indx = 476
    #10;
    addra = 32'd15264;
    dina = {96'd0, 16'd1933, 16'd28980, 16'd60462, 16'd25309, 16'd50839, 16'd9148, 16'd31566, 16'd24407, 16'd53140, 16'd36656}; // indx = 477
    #10;
    addra = 32'd15296;
    dina = {96'd0, 16'd3601, 16'd57222, 16'd34246, 16'd26252, 16'd29459, 16'd8434, 16'd37185, 16'd14741, 16'd18758, 16'd13460}; // indx = 478
    #10;
    addra = 32'd15328;
    dina = {96'd0, 16'd43485, 16'd52304, 16'd49709, 16'd10751, 16'd10745, 16'd40459, 16'd39029, 16'd29965, 16'd6770, 16'd62072}; // indx = 479
    #10;
    addra = 32'd15360;
    dina = {96'd0, 16'd15587, 16'd40505, 16'd30566, 16'd494, 16'd20448, 16'd54566, 16'd5868, 16'd27714, 16'd21745, 16'd14079}; // indx = 480
    #10;
    addra = 32'd15392;
    dina = {96'd0, 16'd53058, 16'd62464, 16'd369, 16'd4142, 16'd24409, 16'd63843, 16'd54424, 16'd21674, 16'd9843, 16'd10058}; // indx = 481
    #10;
    addra = 32'd15424;
    dina = {96'd0, 16'd52328, 16'd35652, 16'd64040, 16'd28505, 16'd11198, 16'd16025, 16'd15436, 16'd10592, 16'd52109, 16'd64055}; // indx = 482
    #10;
    addra = 32'd15456;
    dina = {96'd0, 16'd30970, 16'd9316, 16'd60609, 16'd33537, 16'd62627, 16'd28414, 16'd33616, 16'd61172, 16'd27503, 16'd65208}; // indx = 483
    #10;
    addra = 32'd15488;
    dina = {96'd0, 16'd31914, 16'd57091, 16'd11329, 16'd29578, 16'd58179, 16'd55979, 16'd47791, 16'd6899, 16'd57033, 16'd53475}; // indx = 484
    #10;
    addra = 32'd15520;
    dina = {96'd0, 16'd3078, 16'd52264, 16'd29156, 16'd16396, 16'd44821, 16'd5301, 16'd8352, 16'd32235, 16'd36824, 16'd4871}; // indx = 485
    #10;
    addra = 32'd15552;
    dina = {96'd0, 16'd43808, 16'd47427, 16'd33398, 16'd53322, 16'd43128, 16'd1479, 16'd5476, 16'd58725, 16'd58517, 16'd36241}; // indx = 486
    #10;
    addra = 32'd15584;
    dina = {96'd0, 16'd31454, 16'd3556, 16'd29847, 16'd34045, 16'd60814, 16'd7142, 16'd55459, 16'd56200, 16'd26878, 16'd17276}; // indx = 487
    #10;
    addra = 32'd15616;
    dina = {96'd0, 16'd46989, 16'd14530, 16'd58569, 16'd16782, 16'd38729, 16'd6486, 16'd41022, 16'd47056, 16'd31174, 16'd14058}; // indx = 488
    #10;
    addra = 32'd15648;
    dina = {96'd0, 16'd19613, 16'd15336, 16'd33536, 16'd32513, 16'd4882, 16'd55141, 16'd1468, 16'd38173, 16'd39352, 16'd47360}; // indx = 489
    #10;
    addra = 32'd15680;
    dina = {96'd0, 16'd16495, 16'd52730, 16'd33666, 16'd34799, 16'd24855, 16'd30983, 16'd24506, 16'd17797, 16'd35182, 16'd52498}; // indx = 490
    #10;
    addra = 32'd15712;
    dina = {96'd0, 16'd52331, 16'd55865, 16'd60203, 16'd8306, 16'd8338, 16'd13144, 16'd24540, 16'd59930, 16'd46179, 16'd9158}; // indx = 491
    #10;
    addra = 32'd15744;
    dina = {96'd0, 16'd26920, 16'd39196, 16'd52944, 16'd64346, 16'd11673, 16'd57514, 16'd26436, 16'd1578, 16'd33093, 16'd46813}; // indx = 492
    #10;
    addra = 32'd15776;
    dina = {96'd0, 16'd60013, 16'd4277, 16'd27762, 16'd484, 16'd22534, 16'd65028, 16'd35089, 16'd9801, 16'd23376, 16'd40935}; // indx = 493
    #10;
    addra = 32'd15808;
    dina = {96'd0, 16'd47980, 16'd46089, 16'd62934, 16'd50892, 16'd1016, 16'd16077, 16'd16231, 16'd60700, 16'd38467, 16'd51135}; // indx = 494
    #10;
    addra = 32'd15840;
    dina = {96'd0, 16'd44457, 16'd52648, 16'd4744, 16'd61952, 16'd5112, 16'd46820, 16'd59322, 16'd37569, 16'd18675, 16'd13436}; // indx = 495
    #10;
    addra = 32'd15872;
    dina = {96'd0, 16'd55484, 16'd31837, 16'd59915, 16'd33993, 16'd60720, 16'd44790, 16'd5791, 16'd52316, 16'd16507, 16'd23076}; // indx = 496
    #10;
    addra = 32'd15904;
    dina = {96'd0, 16'd31048, 16'd51930, 16'd62374, 16'd46936, 16'd7153, 16'd14608, 16'd63314, 16'd31702, 16'd7747, 16'd53481}; // indx = 497
    #10;
    addra = 32'd15936;
    dina = {96'd0, 16'd56916, 16'd12366, 16'd25142, 16'd65037, 16'd10981, 16'd57067, 16'd11063, 16'd41278, 16'd63728, 16'd34229}; // indx = 498
    #10;
    addra = 32'd15968;
    dina = {96'd0, 16'd52446, 16'd23848, 16'd18950, 16'd38039, 16'd65080, 16'd21682, 16'd11124, 16'd43412, 16'd56752, 16'd11434}; // indx = 499
    #10;
    addra = 32'd16000;
    dina = {96'd0, 16'd22270, 16'd63621, 16'd35407, 16'd6515, 16'd11247, 16'd46830, 16'd172, 16'd32157, 16'd13870, 16'd56469}; // indx = 500
    #10;
    addra = 32'd16032;
    dina = {96'd0, 16'd64034, 16'd58122, 16'd9916, 16'd26838, 16'd45016, 16'd13078, 16'd62030, 16'd43391, 16'd7395, 16'd20344}; // indx = 501
    #10;
    addra = 32'd16064;
    dina = {96'd0, 16'd61011, 16'd36918, 16'd8067, 16'd58765, 16'd21164, 16'd9900, 16'd4688, 16'd5344, 16'd29610, 16'd58842}; // indx = 502
    #10;
    addra = 32'd16096;
    dina = {96'd0, 16'd23327, 16'd30037, 16'd29654, 16'd21175, 16'd41331, 16'd28848, 16'd38233, 16'd53068, 16'd33319, 16'd45156}; // indx = 503
    #10;
    addra = 32'd16128;
    dina = {96'd0, 16'd46854, 16'd41832, 16'd64774, 16'd16561, 16'd29123, 16'd58631, 16'd47141, 16'd65133, 16'd43147, 16'd15434}; // indx = 504
    #10;
    addra = 32'd16160;
    dina = {96'd0, 16'd48985, 16'd50666, 16'd31268, 16'd6919, 16'd23159, 16'd63998, 16'd60053, 16'd4302, 16'd13080, 16'd44053}; // indx = 505
    #10;
    addra = 32'd16192;
    dina = {96'd0, 16'd65219, 16'd1862, 16'd34880, 16'd19298, 16'd1234, 16'd15753, 16'd158, 16'd4617, 16'd28659, 16'd20703}; // indx = 506
    #10;
    addra = 32'd16224;
    dina = {96'd0, 16'd45024, 16'd31896, 16'd18421, 16'd16808, 16'd49690, 16'd4850, 16'd47821, 16'd15890, 16'd64162, 16'd13461}; // indx = 507
    #10;
    addra = 32'd16256;
    dina = {96'd0, 16'd6331, 16'd8238, 16'd3313, 16'd10897, 16'd40729, 16'd57855, 16'd31431, 16'd38892, 16'd22891, 16'd9813}; // indx = 508
    #10;
    addra = 32'd16288;
    dina = {96'd0, 16'd27699, 16'd12199, 16'd13964, 16'd10780, 16'd47861, 16'd28717, 16'd16967, 16'd36161, 16'd52964, 16'd53232}; // indx = 509
    #10;
    addra = 32'd16320;
    dina = {96'd0, 16'd41760, 16'd65010, 16'd7982, 16'd10504, 16'd26600, 16'd48285, 16'd46677, 16'd12910, 16'd30664, 16'd38577}; // indx = 510
    #10;
    addra = 32'd16352;
    dina = {96'd0, 16'd40158, 16'd9345, 16'd49126, 16'd4657, 16'd44419, 16'd5530, 16'd29350, 16'd40872, 16'd8726, 16'd14816}; // indx = 511
    #10;
    addra = 32'd16384;
    dina = {96'd0, 16'd48792, 16'd4654, 16'd38549, 16'd10003, 16'd59809, 16'd41135, 16'd15478, 16'd23929, 16'd34581, 16'd28169}; // indx = 512
    #10;
    addra = 32'd16416;
    dina = {96'd0, 16'd24992, 16'd50459, 16'd21642, 16'd41453, 16'd11816, 16'd16464, 16'd60145, 16'd18434, 16'd55420, 16'd50329}; // indx = 513
    #10;
    addra = 32'd16448;
    dina = {96'd0, 16'd15638, 16'd42287, 16'd60274, 16'd20381, 16'd57199, 16'd62128, 16'd3237, 16'd61792, 16'd23621, 16'd14907}; // indx = 514
    #10;
    addra = 32'd16480;
    dina = {96'd0, 16'd55889, 16'd5402, 16'd36018, 16'd1552, 16'd1258, 16'd7325, 16'd17647, 16'd40361, 16'd19746, 16'd18925}; // indx = 515
    #10;
    addra = 32'd16512;
    dina = {96'd0, 16'd57469, 16'd10182, 16'd61467, 16'd62473, 16'd4103, 16'd24104, 16'd7252, 16'd33527, 16'd53619, 16'd59780}; // indx = 516
    #10;
    addra = 32'd16544;
    dina = {96'd0, 16'd26978, 16'd39007, 16'd2304, 16'd23, 16'd12047, 16'd57419, 16'd15326, 16'd10653, 16'd21277, 16'd47507}; // indx = 517
    #10;
    addra = 32'd16576;
    dina = {96'd0, 16'd44490, 16'd5017, 16'd5012, 16'd44005, 16'd30123, 16'd36266, 16'd56350, 16'd18355, 16'd31318, 16'd13784}; // indx = 518
    #10;
    addra = 32'd16608;
    dina = {96'd0, 16'd20883, 16'd53424, 16'd60690, 16'd26675, 16'd27347, 16'd40259, 16'd39865, 16'd38881, 16'd46254, 16'd56824}; // indx = 519
    #10;
    addra = 32'd16640;
    dina = {96'd0, 16'd42721, 16'd14838, 16'd36712, 16'd1968, 16'd43909, 16'd40160, 16'd62562, 16'd28483, 16'd22664, 16'd2044}; // indx = 520
    #10;
    addra = 32'd16672;
    dina = {96'd0, 16'd35805, 16'd46369, 16'd38602, 16'd6284, 16'd57018, 16'd39047, 16'd19585, 16'd2528, 16'd21209, 16'd32282}; // indx = 521
    #10;
    addra = 32'd16704;
    dina = {96'd0, 16'd4407, 16'd60392, 16'd55911, 16'd54058, 16'd8711, 16'd25082, 16'd25152, 16'd14247, 16'd39148, 16'd44251}; // indx = 522
    #10;
    addra = 32'd16736;
    dina = {96'd0, 16'd61418, 16'd16681, 16'd59858, 16'd53372, 16'd32642, 16'd20527, 16'd40287, 16'd7825, 16'd20978, 16'd60327}; // indx = 523
    #10;
    addra = 32'd16768;
    dina = {96'd0, 16'd60467, 16'd50934, 16'd40559, 16'd55272, 16'd26184, 16'd50396, 16'd24943, 16'd25794, 16'd8445, 16'd60923}; // indx = 524
    #10;
    addra = 32'd16800;
    dina = {96'd0, 16'd60781, 16'd2671, 16'd42126, 16'd48641, 16'd4479, 16'd56796, 16'd57884, 16'd21128, 16'd5159, 16'd46832}; // indx = 525
    #10;
    addra = 32'd16832;
    dina = {96'd0, 16'd7993, 16'd10174, 16'd30323, 16'd52925, 16'd50624, 16'd8955, 16'd60892, 16'd16511, 16'd12097, 16'd9487}; // indx = 526
    #10;
    addra = 32'd16864;
    dina = {96'd0, 16'd18380, 16'd24151, 16'd37821, 16'd50216, 16'd99, 16'd50191, 16'd2544, 16'd23324, 16'd42823, 16'd54008}; // indx = 527
    #10;
    addra = 32'd16896;
    dina = {96'd0, 16'd56726, 16'd12177, 16'd63750, 16'd6319, 16'd64045, 16'd28779, 16'd21987, 16'd18088, 16'd5559, 16'd50228}; // indx = 528
    #10;
    addra = 32'd16928;
    dina = {96'd0, 16'd4267, 16'd2119, 16'd64896, 16'd46565, 16'd51911, 16'd44014, 16'd45305, 16'd56462, 16'd6664, 16'd33353}; // indx = 529
    #10;
    addra = 32'd16960;
    dina = {96'd0, 16'd1038, 16'd55400, 16'd34791, 16'd65375, 16'd9760, 16'd60868, 16'd48496, 16'd41998, 16'd46585, 16'd30505}; // indx = 530
    #10;
    addra = 32'd16992;
    dina = {96'd0, 16'd51349, 16'd39417, 16'd24773, 16'd56072, 16'd30213, 16'd59561, 16'd53211, 16'd54723, 16'd62297, 16'd25950}; // indx = 531
    #10;
    addra = 32'd17024;
    dina = {96'd0, 16'd25880, 16'd31145, 16'd38264, 16'd27917, 16'd45528, 16'd20597, 16'd39955, 16'd33701, 16'd37523, 16'd43162}; // indx = 532
    #10;
    addra = 32'd17056;
    dina = {96'd0, 16'd22777, 16'd56630, 16'd28003, 16'd38550, 16'd18289, 16'd33640, 16'd2882, 16'd5421, 16'd46030, 16'd9383}; // indx = 533
    #10;
    addra = 32'd17088;
    dina = {96'd0, 16'd49325, 16'd10977, 16'd40062, 16'd24304, 16'd15844, 16'd51575, 16'd31373, 16'd1962, 16'd39175, 16'd44012}; // indx = 534
    #10;
    addra = 32'd17120;
    dina = {96'd0, 16'd47497, 16'd27021, 16'd36532, 16'd50971, 16'd51592, 16'd62492, 16'd39474, 16'd19043, 16'd64688, 16'd20799}; // indx = 535
    #10;
    addra = 32'd17152;
    dina = {96'd0, 16'd2037, 16'd21671, 16'd35347, 16'd36937, 16'd17574, 16'd9714, 16'd9841, 16'd29969, 16'd2412, 16'd5829}; // indx = 536
    #10;
    addra = 32'd17184;
    dina = {96'd0, 16'd50807, 16'd15999, 16'd46878, 16'd58190, 16'd30935, 16'd20067, 16'd47026, 16'd55915, 16'd52181, 16'd21706}; // indx = 537
    #10;
    addra = 32'd17216;
    dina = {96'd0, 16'd54875, 16'd62061, 16'd60346, 16'd3913, 16'd64002, 16'd5921, 16'd44661, 16'd31768, 16'd14984, 16'd31290}; // indx = 538
    #10;
    addra = 32'd17248;
    dina = {96'd0, 16'd29819, 16'd2575, 16'd1070, 16'd1779, 16'd10171, 16'd25823, 16'd13090, 16'd6629, 16'd9997, 16'd26039}; // indx = 539
    #10;
    addra = 32'd17280;
    dina = {96'd0, 16'd22385, 16'd32979, 16'd19962, 16'd38387, 16'd15418, 16'd20583, 16'd28632, 16'd24611, 16'd33708, 16'd63138}; // indx = 540
    #10;
    addra = 32'd17312;
    dina = {96'd0, 16'd42893, 16'd19633, 16'd31355, 16'd75, 16'd9332, 16'd23259, 16'd17434, 16'd28668, 16'd48808, 16'd35690}; // indx = 541
    #10;
    addra = 32'd17344;
    dina = {96'd0, 16'd50131, 16'd16605, 16'd46000, 16'd46988, 16'd62720, 16'd15189, 16'd61127, 16'd52202, 16'd10704, 16'd36139}; // indx = 542
    #10;
    addra = 32'd17376;
    dina = {96'd0, 16'd40725, 16'd8436, 16'd56582, 16'd18922, 16'd2919, 16'd3563, 16'd55783, 16'd19146, 16'd43832, 16'd50655}; // indx = 543
    #10;
    addra = 32'd17408;
    dina = {96'd0, 16'd27829, 16'd46271, 16'd57193, 16'd49024, 16'd21830, 16'd42184, 16'd11874, 16'd50425, 16'd61062, 16'd47696}; // indx = 544
    #10;
    addra = 32'd17440;
    dina = {96'd0, 16'd1887, 16'd4134, 16'd12814, 16'd29675, 16'd51469, 16'd3808, 16'd11149, 16'd58166, 16'd46952, 16'd17398}; // indx = 545
    #10;
    addra = 32'd17472;
    dina = {96'd0, 16'd48842, 16'd31407, 16'd25763, 16'd47902, 16'd30518, 16'd47829, 16'd38250, 16'd41522, 16'd28660, 16'd53959}; // indx = 546
    #10;
    addra = 32'd17504;
    dina = {96'd0, 16'd17627, 16'd21359, 16'd21328, 16'd30882, 16'd32014, 16'd14770, 16'd173, 16'd45685, 16'd53509, 16'd53812}; // indx = 547
    #10;
    addra = 32'd17536;
    dina = {96'd0, 16'd17199, 16'd20083, 16'd20196, 16'd10341, 16'd44749, 16'd17054, 16'd31094, 16'd52088, 16'd36906, 16'd62726}; // indx = 548
    #10;
    addra = 32'd17568;
    dina = {96'd0, 16'd17649, 16'd53490, 16'd28986, 16'd22278, 16'd28940, 16'd15188, 16'd55152, 16'd33174, 16'd35207, 16'd1339}; // indx = 549
    #10;
    addra = 32'd17600;
    dina = {96'd0, 16'd59758, 16'd37923, 16'd35794, 16'd39431, 16'd12128, 16'd45018, 16'd21407, 16'd13859, 16'd62657, 16'd21336}; // indx = 550
    #10;
    addra = 32'd17632;
    dina = {96'd0, 16'd28671, 16'd59650, 16'd9996, 16'd5337, 16'd47575, 16'd50391, 16'd25924, 16'd62811, 16'd60091, 16'd3190}; // indx = 551
    #10;
    addra = 32'd17664;
    dina = {96'd0, 16'd18144, 16'd4259, 16'd18612, 16'd62976, 16'd41716, 16'd21561, 16'd44838, 16'd1495, 16'd58836, 16'd33160}; // indx = 552
    #10;
    addra = 32'd17696;
    dina = {96'd0, 16'd11691, 16'd59515, 16'd50579, 16'd61247, 16'd64109, 16'd62858, 16'd11525, 16'd44504, 16'd17677, 16'd50032}; // indx = 553
    #10;
    addra = 32'd17728;
    dina = {96'd0, 16'd60910, 16'd44053, 16'd27263, 16'd28517, 16'd59105, 16'd45432, 16'd26149, 16'd7753, 16'd30858, 16'd20484}; // indx = 554
    #10;
    addra = 32'd17760;
    dina = {96'd0, 16'd40997, 16'd64910, 16'd62899, 16'd8367, 16'd39644, 16'd1206, 16'd45286, 16'd42908, 16'd43968, 16'd49392}; // indx = 555
    #10;
    addra = 32'd17792;
    dina = {96'd0, 16'd27626, 16'd53877, 16'd49903, 16'd55739, 16'd43301, 16'd5269, 16'd18110, 16'd53423, 16'd14733, 16'd4119}; // indx = 556
    #10;
    addra = 32'd17824;
    dina = {96'd0, 16'd20143, 16'd34934, 16'd52693, 16'd58237, 16'd36116, 16'd56112, 16'd55680, 16'd6775, 16'd20276, 16'd47133}; // indx = 557
    #10;
    addra = 32'd17856;
    dina = {96'd0, 16'd32033, 16'd46551, 16'd50630, 16'd28062, 16'd25952, 16'd50412, 16'd22737, 16'd57293, 16'd6052, 16'd64350}; // indx = 558
    #10;
    addra = 32'd17888;
    dina = {96'd0, 16'd22379, 16'd35880, 16'd2647, 16'd37985, 16'd43934, 16'd2143, 16'd61647, 16'd44661, 16'd34380, 16'd21288}; // indx = 559
    #10;
    addra = 32'd17920;
    dina = {96'd0, 16'd28148, 16'd15897, 16'd7093, 16'd5736, 16'd40921, 16'd4742, 16'd7996, 16'd9026, 16'd26870, 16'd1742}; // indx = 560
    #10;
    addra = 32'd17952;
    dina = {96'd0, 16'd20824, 16'd46657, 16'd61315, 16'd4170, 16'd44877, 16'd37239, 16'd33022, 16'd48891, 16'd45004, 16'd15917}; // indx = 561
    #10;
    addra = 32'd17984;
    dina = {96'd0, 16'd1862, 16'd24508, 16'd41353, 16'd57268, 16'd28095, 16'd41541, 16'd21468, 16'd3872, 16'd42348, 16'd5074}; // indx = 562
    #10;
    addra = 32'd18016;
    dina = {96'd0, 16'd23994, 16'd52219, 16'd17664, 16'd10657, 16'd8005, 16'd22078, 16'd22006, 16'd5776, 16'd6026, 16'd35157}; // indx = 563
    #10;
    addra = 32'd18048;
    dina = {96'd0, 16'd61432, 16'd39406, 16'd60844, 16'd13947, 16'd47389, 16'd15716, 16'd24700, 16'd32732, 16'd54262, 16'd412}; // indx = 564
    #10;
    addra = 32'd18080;
    dina = {96'd0, 16'd21609, 16'd34012, 16'd8249, 16'd28658, 16'd39394, 16'd26175, 16'd45775, 16'd43925, 16'd56632, 16'd50037}; // indx = 565
    #10;
    addra = 32'd18112;
    dina = {96'd0, 16'd59437, 16'd30717, 16'd64356, 16'd57892, 16'd45019, 16'd8718, 16'd30658, 16'd29440, 16'd13955, 16'd48248}; // indx = 566
    #10;
    addra = 32'd18144;
    dina = {96'd0, 16'd42824, 16'd19934, 16'd38793, 16'd45081, 16'd10176, 16'd16398, 16'd31651, 16'd39566, 16'd34264, 16'd44464}; // indx = 567
    #10;
    addra = 32'd18176;
    dina = {96'd0, 16'd32547, 16'd25394, 16'd6803, 16'd32988, 16'd42895, 16'd64669, 16'd38302, 16'd60090, 16'd19680, 16'd56032}; // indx = 568
    #10;
    addra = 32'd18208;
    dina = {96'd0, 16'd24757, 16'd41373, 16'd59490, 16'd55237, 16'd50197, 16'd49017, 16'd53574, 16'd17819, 16'd51592, 16'd10137}; // indx = 569
    #10;
    addra = 32'd18240;
    dina = {96'd0, 16'd3970, 16'd8519, 16'd26236, 16'd40234, 16'd32004, 16'd5283, 16'd63619, 16'd31895, 16'd24379, 16'd29869}; // indx = 570
    #10;
    addra = 32'd18272;
    dina = {96'd0, 16'd56444, 16'd4292, 16'd41167, 16'd50806, 16'd3981, 16'd52919, 16'd57735, 16'd4130, 16'd45898, 16'd62936}; // indx = 571
    #10;
    addra = 32'd18304;
    dina = {96'd0, 16'd11280, 16'd53714, 16'd63253, 16'd59984, 16'd15993, 16'd35398, 16'd40425, 16'd42214, 16'd52651, 16'd28625}; // indx = 572
    #10;
    addra = 32'd18336;
    dina = {96'd0, 16'd5540, 16'd9505, 16'd40986, 16'd23072, 16'd13918, 16'd64480, 16'd43677, 16'd39659, 16'd1585, 16'd65342}; // indx = 573
    #10;
    addra = 32'd18368;
    dina = {96'd0, 16'd33406, 16'd45921, 16'd26209, 16'd40243, 16'd1471, 16'd55151, 16'd51158, 16'd8798, 16'd14227, 16'd50631}; // indx = 574
    #10;
    addra = 32'd18400;
    dina = {96'd0, 16'd42964, 16'd34928, 16'd5266, 16'd56606, 16'd1897, 16'd45733, 16'd56452, 16'd14564, 16'd52768, 16'd35941}; // indx = 575
    #10;
    addra = 32'd18432;
    dina = {96'd0, 16'd6335, 16'd59746, 16'd45552, 16'd23636, 16'd27757, 16'd61955, 16'd15434, 16'd41244, 16'd44493, 16'd51350}; // indx = 576
    #10;
    addra = 32'd18464;
    dina = {96'd0, 16'd7981, 16'd10175, 16'd36676, 16'd60835, 16'd40181, 16'd15827, 16'd34793, 16'd36474, 16'd9768, 16'd54573}; // indx = 577
    #10;
    addra = 32'd18496;
    dina = {96'd0, 16'd54030, 16'd34442, 16'd36856, 16'd52339, 16'd51468, 16'd21629, 16'd9928, 16'd2730, 16'd40921, 16'd17455}; // indx = 578
    #10;
    addra = 32'd18528;
    dina = {96'd0, 16'd59312, 16'd58286, 16'd5176, 16'd12907, 16'd32066, 16'd40911, 16'd64490, 16'd36573, 16'd30417, 16'd28640}; // indx = 579
    #10;
    addra = 32'd18560;
    dina = {96'd0, 16'd17640, 16'd12030, 16'd51633, 16'd35568, 16'd2456, 16'd2926, 16'd51218, 16'd32193, 16'd2235, 16'd30780}; // indx = 580
    #10;
    addra = 32'd18592;
    dina = {96'd0, 16'd11610, 16'd53960, 16'd56688, 16'd22219, 16'd3486, 16'd4105, 16'd22568, 16'd62129, 16'd48351, 16'd28985}; // indx = 581
    #10;
    addra = 32'd18624;
    dina = {96'd0, 16'd10616, 16'd14481, 16'd46840, 16'd62046, 16'd65310, 16'd33079, 16'd56256, 16'd64343, 16'd53218, 16'd11520}; // indx = 582
    #10;
    addra = 32'd18656;
    dina = {96'd0, 16'd56313, 16'd51310, 16'd25648, 16'd60537, 16'd38898, 16'd33909, 16'd53680, 16'd38840, 16'd43601, 16'd51195}; // indx = 583
    #10;
    addra = 32'd18688;
    dina = {96'd0, 16'd27742, 16'd34134, 16'd54027, 16'd2382, 16'd5467, 16'd5724, 16'd17775, 16'd40617, 16'd59926, 16'd61928}; // indx = 584
    #10;
    addra = 32'd18720;
    dina = {96'd0, 16'd45481, 16'd32876, 16'd10023, 16'd746, 16'd1451, 16'd49110, 16'd25285, 16'd7327, 16'd57940, 16'd65031}; // indx = 585
    #10;
    addra = 32'd18752;
    dina = {96'd0, 16'd19156, 16'd45201, 16'd54220, 16'd57447, 16'd27663, 16'd11460, 16'd39820, 16'd34726, 16'd31780, 16'd10537}; // indx = 586
    #10;
    addra = 32'd18784;
    dina = {96'd0, 16'd17404, 16'd59547, 16'd18485, 16'd55663, 16'd3387, 16'd21382, 16'd63604, 16'd55121, 16'd36508, 16'd34693}; // indx = 587
    #10;
    addra = 32'd18816;
    dina = {96'd0, 16'd26830, 16'd53473, 16'd3628, 16'd19009, 16'd57626, 16'd59784, 16'd33293, 16'd168, 16'd58831, 16'd35450}; // indx = 588
    #10;
    addra = 32'd18848;
    dina = {96'd0, 16'd44444, 16'd49825, 16'd10365, 16'd11140, 16'd30397, 16'd4704, 16'd49852, 16'd29246, 16'd46760, 16'd2439}; // indx = 589
    #10;
    addra = 32'd18880;
    dina = {96'd0, 16'd65513, 16'd23678, 16'd16361, 16'd57856, 16'd2222, 16'd6984, 16'd26748, 16'd7864, 16'd41681, 16'd46799}; // indx = 590
    #10;
    addra = 32'd18912;
    dina = {96'd0, 16'd8345, 16'd15251, 16'd8775, 16'd53401, 16'd16057, 16'd16354, 16'd59596, 16'd37015, 16'd57048, 16'd56897}; // indx = 591
    #10;
    addra = 32'd18944;
    dina = {96'd0, 16'd35954, 16'd7112, 16'd43157, 16'd42000, 16'd45659, 16'd23861, 16'd58614, 16'd21516, 16'd15346, 16'd26915}; // indx = 592
    #10;
    addra = 32'd18976;
    dina = {96'd0, 16'd24748, 16'd40163, 16'd21498, 16'd23166, 16'd51632, 16'd57082, 16'd51852, 16'd10666, 16'd63500, 16'd20138}; // indx = 593
    #10;
    addra = 32'd19008;
    dina = {96'd0, 16'd39896, 16'd24867, 16'd29038, 16'd16616, 16'd2195, 16'd59178, 16'd4489, 16'd21290, 16'd50956, 16'd56383}; // indx = 594
    #10;
    addra = 32'd19040;
    dina = {96'd0, 16'd32325, 16'd58598, 16'd31002, 16'd63260, 16'd28318, 16'd41253, 16'd50367, 16'd50251, 16'd54163, 16'd64931}; // indx = 595
    #10;
    addra = 32'd19072;
    dina = {96'd0, 16'd53855, 16'd29011, 16'd19329, 16'd17490, 16'd40152, 16'd9709, 16'd1363, 16'd48867, 16'd8220, 16'd65087}; // indx = 596
    #10;
    addra = 32'd19104;
    dina = {96'd0, 16'd5976, 16'd3292, 16'd45972, 16'd60698, 16'd15685, 16'd48373, 16'd43114, 16'd51650, 16'd51190, 16'd1517}; // indx = 597
    #10;
    addra = 32'd19136;
    dina = {96'd0, 16'd1464, 16'd7931, 16'd61870, 16'd31764, 16'd61830, 16'd61533, 16'd29108, 16'd18362, 16'd56364, 16'd61314}; // indx = 598
    #10;
    addra = 32'd19168;
    dina = {96'd0, 16'd21904, 16'd44883, 16'd13715, 16'd13165, 16'd15511, 16'd54137, 16'd24400, 16'd989, 16'd32982, 16'd2644}; // indx = 599
    #10;
    addra = 32'd19200;
    dina = {96'd0, 16'd10198, 16'd12442, 16'd55497, 16'd45751, 16'd1613, 16'd28956, 16'd53129, 16'd42971, 16'd29078, 16'd36623}; // indx = 600
    #10;
    addra = 32'd19232;
    dina = {96'd0, 16'd59749, 16'd16202, 16'd31500, 16'd23392, 16'd60237, 16'd10936, 16'd20479, 16'd6458, 16'd10100, 16'd36832}; // indx = 601
    #10;
    addra = 32'd19264;
    dina = {96'd0, 16'd18617, 16'd52325, 16'd14593, 16'd60776, 16'd8729, 16'd49360, 16'd18430, 16'd22018, 16'd57740, 16'd19822}; // indx = 602
    #10;
    addra = 32'd19296;
    dina = {96'd0, 16'd21215, 16'd65525, 16'd21268, 16'd51665, 16'd25759, 16'd41921, 16'd17311, 16'd38445, 16'd19189, 16'd19864}; // indx = 603
    #10;
    addra = 32'd19328;
    dina = {96'd0, 16'd34037, 16'd26593, 16'd52653, 16'd20560, 16'd17972, 16'd42870, 16'd57597, 16'd22466, 16'd65055, 16'd16906}; // indx = 604
    #10;
    addra = 32'd19360;
    dina = {96'd0, 16'd23348, 16'd11488, 16'd58006, 16'd5709, 16'd4944, 16'd872, 16'd44477, 16'd1383, 16'd23727, 16'd18730}; // indx = 605
    #10;
    addra = 32'd19392;
    dina = {96'd0, 16'd56767, 16'd63883, 16'd5583, 16'd48464, 16'd2154, 16'd11375, 16'd4973, 16'd13716, 16'd54516, 16'd16076}; // indx = 606
    #10;
    addra = 32'd19424;
    dina = {96'd0, 16'd27542, 16'd37495, 16'd30733, 16'd21066, 16'd31805, 16'd54091, 16'd8589, 16'd52491, 16'd58698, 16'd38051}; // indx = 607
    #10;
    addra = 32'd19456;
    dina = {96'd0, 16'd26557, 16'd54691, 16'd61774, 16'd64768, 16'd16612, 16'd40621, 16'd40301, 16'd52446, 16'd55122, 16'd48331}; // indx = 608
    #10;
    addra = 32'd19488;
    dina = {96'd0, 16'd39833, 16'd52536, 16'd12862, 16'd47949, 16'd13205, 16'd29094, 16'd25541, 16'd2137, 16'd41504, 16'd55639}; // indx = 609
    #10;
    addra = 32'd19520;
    dina = {96'd0, 16'd51697, 16'd29476, 16'd21952, 16'd64334, 16'd5946, 16'd841, 16'd6382, 16'd28888, 16'd3520, 16'd6474}; // indx = 610
    #10;
    addra = 32'd19552;
    dina = {96'd0, 16'd26115, 16'd24247, 16'd59819, 16'd24937, 16'd55947, 16'd30855, 16'd43343, 16'd30855, 16'd56580, 16'd39789}; // indx = 611
    #10;
    addra = 32'd19584;
    dina = {96'd0, 16'd40461, 16'd62474, 16'd63358, 16'd65226, 16'd26206, 16'd5058, 16'd64932, 16'd13859, 16'd8396, 16'd48931}; // indx = 612
    #10;
    addra = 32'd19616;
    dina = {96'd0, 16'd38491, 16'd7129, 16'd24705, 16'd47257, 16'd60143, 16'd51655, 16'd54951, 16'd52680, 16'd21753, 16'd36010}; // indx = 613
    #10;
    addra = 32'd19648;
    dina = {96'd0, 16'd64330, 16'd15533, 16'd45668, 16'd6519, 16'd49053, 16'd17357, 16'd11247, 16'd32229, 16'd1762, 16'd5906}; // indx = 614
    #10;
    addra = 32'd19680;
    dina = {96'd0, 16'd53920, 16'd963, 16'd59322, 16'd19312, 16'd33122, 16'd58958, 16'd42761, 16'd27273, 16'd22979, 16'd29533}; // indx = 615
    #10;
    addra = 32'd19712;
    dina = {96'd0, 16'd18784, 16'd46172, 16'd55278, 16'd31679, 16'd7856, 16'd14883, 16'd41088, 16'd62235, 16'd12017, 16'd51278}; // indx = 616
    #10;
    addra = 32'd19744;
    dina = {96'd0, 16'd22761, 16'd16890, 16'd34763, 16'd48616, 16'd50568, 16'd18165, 16'd38023, 16'd65482, 16'd54611, 16'd13473}; // indx = 617
    #10;
    addra = 32'd19776;
    dina = {96'd0, 16'd24562, 16'd47900, 16'd10422, 16'd41205, 16'd8233, 16'd7423, 16'd40865, 16'd28117, 16'd52157, 16'd57798}; // indx = 618
    #10;
    addra = 32'd19808;
    dina = {96'd0, 16'd7464, 16'd22576, 16'd401, 16'd21082, 16'd56951, 16'd34579, 16'd31373, 16'd7016, 16'd22440, 16'd1910}; // indx = 619
    #10;
    addra = 32'd19840;
    dina = {96'd0, 16'd49110, 16'd36200, 16'd11694, 16'd26267, 16'd21901, 16'd62150, 16'd59863, 16'd24183, 16'd39953, 16'd19246}; // indx = 620
    #10;
    addra = 32'd19872;
    dina = {96'd0, 16'd55353, 16'd2853, 16'd43738, 16'd4424, 16'd54224, 16'd54366, 16'd14533, 16'd13030, 16'd11914, 16'd24605}; // indx = 621
    #10;
    addra = 32'd19904;
    dina = {96'd0, 16'd35328, 16'd4751, 16'd55291, 16'd65525, 16'd12708, 16'd4523, 16'd39563, 16'd16480, 16'd51574, 16'd31650}; // indx = 622
    #10;
    addra = 32'd19936;
    dina = {96'd0, 16'd1362, 16'd10926, 16'd51052, 16'd19026, 16'd3103, 16'd11510, 16'd55745, 16'd23531, 16'd11204, 16'd41867}; // indx = 623
    #10;
    addra = 32'd19968;
    dina = {96'd0, 16'd30660, 16'd42340, 16'd12377, 16'd51376, 16'd17913, 16'd14090, 16'd11458, 16'd19263, 16'd53795, 16'd61211}; // indx = 624
    #10;
    addra = 32'd20000;
    dina = {96'd0, 16'd15998, 16'd45336, 16'd5769, 16'd5555, 16'd3176, 16'd55841, 16'd36656, 16'd52992, 16'd51924, 16'd6728}; // indx = 625
    #10;
    addra = 32'd20032;
    dina = {96'd0, 16'd16921, 16'd53015, 16'd31083, 16'd51408, 16'd15225, 16'd31073, 16'd13566, 16'd50720, 16'd14191, 16'd12731}; // indx = 626
    #10;
    addra = 32'd20064;
    dina = {96'd0, 16'd58967, 16'd39388, 16'd53960, 16'd14111, 16'd6110, 16'd3935, 16'd38161, 16'd29074, 16'd40170, 16'd9009}; // indx = 627
    #10;
    addra = 32'd20096;
    dina = {96'd0, 16'd8677, 16'd27746, 16'd22034, 16'd40334, 16'd37659, 16'd42164, 16'd53830, 16'd23681, 16'd31154, 16'd23171}; // indx = 628
    #10;
    addra = 32'd20128;
    dina = {96'd0, 16'd60608, 16'd7421, 16'd51650, 16'd21124, 16'd23484, 16'd2467, 16'd62151, 16'd19892, 16'd38801, 16'd16437}; // indx = 629
    #10;
    addra = 32'd20160;
    dina = {96'd0, 16'd49861, 16'd2676, 16'd39965, 16'd38368, 16'd60174, 16'd56054, 16'd55380, 16'd22933, 16'd25822, 16'd53527}; // indx = 630
    #10;
    addra = 32'd20192;
    dina = {96'd0, 16'd16180, 16'd41123, 16'd38952, 16'd42935, 16'd36326, 16'd22382, 16'd17487, 16'd24010, 16'd12748, 16'd19526}; // indx = 631
    #10;
    addra = 32'd20224;
    dina = {96'd0, 16'd56417, 16'd24199, 16'd171, 16'd12349, 16'd53612, 16'd60489, 16'd62086, 16'd34285, 16'd10621, 16'd4626}; // indx = 632
    #10;
    addra = 32'd20256;
    dina = {96'd0, 16'd2545, 16'd48074, 16'd28178, 16'd61664, 16'd61578, 16'd45328, 16'd26821, 16'd23690, 16'd11705, 16'd23418}; // indx = 633
    #10;
    addra = 32'd20288;
    dina = {96'd0, 16'd52229, 16'd52544, 16'd34762, 16'd18754, 16'd18100, 16'd5496, 16'd12057, 16'd10580, 16'd11776, 16'd53836}; // indx = 634
    #10;
    addra = 32'd20320;
    dina = {96'd0, 16'd64864, 16'd50342, 16'd12742, 16'd47056, 16'd17853, 16'd49461, 16'd16859, 16'd20354, 16'd21261, 16'd19107}; // indx = 635
    #10;
    addra = 32'd20352;
    dina = {96'd0, 16'd19076, 16'd30416, 16'd12035, 16'd49430, 16'd38807, 16'd51847, 16'd49850, 16'd38227, 16'd7316, 16'd53262}; // indx = 636
    #10;
    addra = 32'd20384;
    dina = {96'd0, 16'd36749, 16'd10526, 16'd9721, 16'd41363, 16'd56214, 16'd36064, 16'd51058, 16'd15522, 16'd20511, 16'd52746}; // indx = 637
    #10;
    addra = 32'd20416;
    dina = {96'd0, 16'd5411, 16'd49343, 16'd19428, 16'd44664, 16'd56141, 16'd27532, 16'd7878, 16'd3822, 16'd28594, 16'd14547}; // indx = 638
    #10;
    addra = 32'd20448;
    dina = {96'd0, 16'd13695, 16'd40242, 16'd24026, 16'd20615, 16'd9387, 16'd1255, 16'd64832, 16'd36129, 16'd29369, 16'd44111}; // indx = 639
    #10;
    addra = 32'd20480;
    dina = {96'd0, 16'd53755, 16'd24992, 16'd43121, 16'd9480, 16'd33141, 16'd7126, 16'd31155, 16'd33906, 16'd44250, 16'd9246}; // indx = 640
    #10;
    addra = 32'd20512;
    dina = {96'd0, 16'd26555, 16'd32384, 16'd18490, 16'd38598, 16'd43788, 16'd17412, 16'd33588, 16'd34387, 16'd5213, 16'd64909}; // indx = 641
    #10;
    addra = 32'd20544;
    dina = {96'd0, 16'd51639, 16'd49239, 16'd34049, 16'd21543, 16'd52826, 16'd63488, 16'd38818, 16'd4184, 16'd42214, 16'd24872}; // indx = 642
    #10;
    addra = 32'd20576;
    dina = {96'd0, 16'd47467, 16'd48714, 16'd53856, 16'd57098, 16'd17895, 16'd54581, 16'd8653, 16'd54430, 16'd19063, 16'd44482}; // indx = 643
    #10;
    addra = 32'd20608;
    dina = {96'd0, 16'd489, 16'd41003, 16'd36815, 16'd7841, 16'd40073, 16'd33073, 16'd846, 16'd60502, 16'd9593, 16'd44436}; // indx = 644
    #10;
    addra = 32'd20640;
    dina = {96'd0, 16'd61134, 16'd44747, 16'd58420, 16'd41246, 16'd2795, 16'd4450, 16'd24005, 16'd63867, 16'd38370, 16'd58975}; // indx = 645
    #10;
    addra = 32'd20672;
    dina = {96'd0, 16'd22396, 16'd16910, 16'd49781, 16'd42657, 16'd3970, 16'd2288, 16'd29042, 16'd6966, 16'd4598, 16'd34553}; // indx = 646
    #10;
    addra = 32'd20704;
    dina = {96'd0, 16'd30203, 16'd41067, 16'd43927, 16'd50907, 16'd57590, 16'd20085, 16'd32584, 16'd36420, 16'd32944, 16'd59890}; // indx = 647
    #10;
    addra = 32'd20736;
    dina = {96'd0, 16'd63066, 16'd11277, 16'd20554, 16'd35646, 16'd49, 16'd17557, 16'd59893, 16'd56221, 16'd50219, 16'd57209}; // indx = 648
    #10;
    addra = 32'd20768;
    dina = {96'd0, 16'd56594, 16'd61802, 16'd17650, 16'd13568, 16'd8747, 16'd19811, 16'd40518, 16'd45060, 16'd56681, 16'd49620}; // indx = 649
    #10;
    addra = 32'd20800;
    dina = {96'd0, 16'd50144, 16'd25143, 16'd27406, 16'd51049, 16'd43130, 16'd46329, 16'd8906, 16'd6910, 16'd17655, 16'd53774}; // indx = 650
    #10;
    addra = 32'd20832;
    dina = {96'd0, 16'd10160, 16'd35416, 16'd47980, 16'd48868, 16'd1144, 16'd60619, 16'd47268, 16'd33861, 16'd45949, 16'd60708}; // indx = 651
    #10;
    addra = 32'd20864;
    dina = {96'd0, 16'd23231, 16'd16088, 16'd836, 16'd28045, 16'd23428, 16'd43612, 16'd17859, 16'd44312, 16'd28358, 16'd10433}; // indx = 652
    #10;
    addra = 32'd20896;
    dina = {96'd0, 16'd11205, 16'd52408, 16'd59400, 16'd42187, 16'd42123, 16'd39807, 16'd48057, 16'd62542, 16'd33732, 16'd6095}; // indx = 653
    #10;
    addra = 32'd20928;
    dina = {96'd0, 16'd34500, 16'd60843, 16'd30135, 16'd38980, 16'd64212, 16'd21913, 16'd34510, 16'd840, 16'd36264, 16'd19842}; // indx = 654
    #10;
    addra = 32'd20960;
    dina = {96'd0, 16'd38692, 16'd36351, 16'd32350, 16'd27145, 16'd32163, 16'd60388, 16'd45135, 16'd50905, 16'd49412, 16'd62428}; // indx = 655
    #10;
    addra = 32'd20992;
    dina = {96'd0, 16'd41731, 16'd57163, 16'd11843, 16'd24923, 16'd14320, 16'd34256, 16'd31638, 16'd29667, 16'd18500, 16'd52764}; // indx = 656
    #10;
    addra = 32'd21024;
    dina = {96'd0, 16'd49098, 16'd2833, 16'd59418, 16'd47678, 16'd58840, 16'd16248, 16'd52851, 16'd30810, 16'd17559, 16'd6914}; // indx = 657
    #10;
    addra = 32'd21056;
    dina = {96'd0, 16'd63812, 16'd9896, 16'd57352, 16'd61582, 16'd54818, 16'd33847, 16'd46735, 16'd57152, 16'd64533, 16'd48272}; // indx = 658
    #10;
    addra = 32'd21088;
    dina = {96'd0, 16'd22781, 16'd40303, 16'd21630, 16'd49734, 16'd12980, 16'd32694, 16'd26475, 16'd60483, 16'd51308, 16'd5038}; // indx = 659
    #10;
    addra = 32'd21120;
    dina = {96'd0, 16'd37221, 16'd23274, 16'd26985, 16'd58713, 16'd51536, 16'd34794, 16'd18598, 16'd15564, 16'd30852, 16'd65516}; // indx = 660
    #10;
    addra = 32'd21152;
    dina = {96'd0, 16'd40841, 16'd24136, 16'd30598, 16'd32859, 16'd36108, 16'd41028, 16'd48941, 16'd28158, 16'd45016, 16'd47825}; // indx = 661
    #10;
    addra = 32'd21184;
    dina = {96'd0, 16'd6454, 16'd58833, 16'd50833, 16'd19388, 16'd3698, 16'd62827, 16'd33458, 16'd6918, 16'd64646, 16'd30126}; // indx = 662
    #10;
    addra = 32'd21216;
    dina = {96'd0, 16'd27024, 16'd50042, 16'd6123, 16'd47591, 16'd24367, 16'd14194, 16'd45051, 16'd27697, 16'd45361, 16'd51048}; // indx = 663
    #10;
    addra = 32'd21248;
    dina = {96'd0, 16'd34418, 16'd22871, 16'd29731, 16'd30636, 16'd38193, 16'd37361, 16'd14231, 16'd20878, 16'd32737, 16'd45953}; // indx = 664
    #10;
    addra = 32'd21280;
    dina = {96'd0, 16'd59379, 16'd57724, 16'd28311, 16'd31995, 16'd53632, 16'd9243, 16'd9738, 16'd61681, 16'd2288, 16'd9242}; // indx = 665
    #10;
    addra = 32'd21312;
    dina = {96'd0, 16'd8939, 16'd38061, 16'd21521, 16'd34836, 16'd4404, 16'd55944, 16'd20056, 16'd34944, 16'd34189, 16'd34736}; // indx = 666
    #10;
    addra = 32'd21344;
    dina = {96'd0, 16'd64490, 16'd57099, 16'd45893, 16'd22150, 16'd45096, 16'd45485, 16'd44687, 16'd38540, 16'd19673, 16'd52123}; // indx = 667
    #10;
    addra = 32'd21376;
    dina = {96'd0, 16'd21872, 16'd62812, 16'd18722, 16'd27535, 16'd39881, 16'd17044, 16'd21290, 16'd50446, 16'd37852, 16'd30668}; // indx = 668
    #10;
    addra = 32'd21408;
    dina = {96'd0, 16'd1647, 16'd37092, 16'd19075, 16'd1109, 16'd61283, 16'd598, 16'd2045, 16'd42790, 16'd17707, 16'd28282}; // indx = 669
    #10;
    addra = 32'd21440;
    dina = {96'd0, 16'd61034, 16'd46399, 16'd49053, 16'd18540, 16'd65471, 16'd33880, 16'd26696, 16'd5143, 16'd49544, 16'd13029}; // indx = 670
    #10;
    addra = 32'd21472;
    dina = {96'd0, 16'd30578, 16'd30702, 16'd62761, 16'd38380, 16'd54980, 16'd4095, 16'd63165, 16'd33952, 16'd18216, 16'd44220}; // indx = 671
    #10;
    addra = 32'd21504;
    dina = {96'd0, 16'd37211, 16'd5716, 16'd35580, 16'd9078, 16'd34218, 16'd12001, 16'd62565, 16'd13835, 16'd21465, 16'd4445}; // indx = 672
    #10;
    addra = 32'd21536;
    dina = {96'd0, 16'd42380, 16'd46208, 16'd13366, 16'd57076, 16'd698, 16'd14705, 16'd48207, 16'd59845, 16'd25861, 16'd12851}; // indx = 673
    #10;
    addra = 32'd21568;
    dina = {96'd0, 16'd57111, 16'd49503, 16'd12466, 16'd19178, 16'd63622, 16'd35395, 16'd42761, 16'd56236, 16'd63424, 16'd9211}; // indx = 674
    #10;
    addra = 32'd21600;
    dina = {96'd0, 16'd45284, 16'd3062, 16'd61153, 16'd50556, 16'd14196, 16'd28215, 16'd36922, 16'd11073, 16'd40249, 16'd34144}; // indx = 675
    #10;
    addra = 32'd21632;
    dina = {96'd0, 16'd9234, 16'd2587, 16'd44071, 16'd53995, 16'd41707, 16'd47825, 16'd48520, 16'd50394, 16'd31551, 16'd33780}; // indx = 676
    #10;
    addra = 32'd21664;
    dina = {96'd0, 16'd33698, 16'd41219, 16'd27255, 16'd53477, 16'd15626, 16'd20134, 16'd6357, 16'd48138, 16'd375, 16'd56607}; // indx = 677
    #10;
    addra = 32'd21696;
    dina = {96'd0, 16'd15307, 16'd23844, 16'd40774, 16'd45966, 16'd6709, 16'd13904, 16'd27460, 16'd62774, 16'd16812, 16'd16863}; // indx = 678
    #10;
    addra = 32'd21728;
    dina = {96'd0, 16'd19941, 16'd63673, 16'd53536, 16'd6530, 16'd17584, 16'd61602, 16'd47492, 16'd1593, 16'd9172, 16'd21428}; // indx = 679
    #10;
    addra = 32'd21760;
    dina = {96'd0, 16'd9536, 16'd57266, 16'd34465, 16'd16705, 16'd3929, 16'd31721, 16'd60956, 16'd25052, 16'd58144, 16'd47055}; // indx = 680
    #10;
    addra = 32'd21792;
    dina = {96'd0, 16'd48348, 16'd23815, 16'd50281, 16'd31330, 16'd28232, 16'd54279, 16'd55528, 16'd43082, 16'd34643, 16'd38003}; // indx = 681
    #10;
    addra = 32'd21824;
    dina = {96'd0, 16'd50812, 16'd55241, 16'd9007, 16'd25930, 16'd62941, 16'd11095, 16'd45078, 16'd54805, 16'd589, 16'd27145}; // indx = 682
    #10;
    addra = 32'd21856;
    dina = {96'd0, 16'd62919, 16'd43040, 16'd62537, 16'd32032, 16'd14325, 16'd15472, 16'd40416, 16'd13634, 16'd25209, 16'd12634}; // indx = 683
    #10;
    addra = 32'd21888;
    dina = {96'd0, 16'd21941, 16'd48190, 16'd50032, 16'd6527, 16'd64163, 16'd31510, 16'd4374, 16'd39724, 16'd37054, 16'd38101}; // indx = 684
    #10;
    addra = 32'd21920;
    dina = {96'd0, 16'd60992, 16'd14334, 16'd42225, 16'd26767, 16'd24441, 16'd19536, 16'd28405, 16'd53767, 16'd51314, 16'd51385}; // indx = 685
    #10;
    addra = 32'd21952;
    dina = {96'd0, 16'd41221, 16'd35273, 16'd22486, 16'd62675, 16'd18166, 16'd58158, 16'd23525, 16'd8700, 16'd54980, 16'd51885}; // indx = 686
    #10;
    addra = 32'd21984;
    dina = {96'd0, 16'd31789, 16'd48786, 16'd49810, 16'd42131, 16'd11502, 16'd64001, 16'd15487, 16'd35343, 16'd37343, 16'd46188}; // indx = 687
    #10;
    addra = 32'd22016;
    dina = {96'd0, 16'd11387, 16'd60737, 16'd9795, 16'd14860, 16'd14755, 16'd24712, 16'd36357, 16'd54497, 16'd43066, 16'd58821}; // indx = 688
    #10;
    addra = 32'd22048;
    dina = {96'd0, 16'd59302, 16'd43671, 16'd41724, 16'd35536, 16'd27899, 16'd8617, 16'd39636, 16'd37215, 16'd61570, 16'd53041}; // indx = 689
    #10;
    addra = 32'd22080;
    dina = {96'd0, 16'd57290, 16'd10913, 16'd16335, 16'd11247, 16'd64289, 16'd46738, 16'd45702, 16'd37571, 16'd24100, 16'd22882}; // indx = 690
    #10;
    addra = 32'd22112;
    dina = {96'd0, 16'd48145, 16'd33795, 16'd5861, 16'd59457, 16'd39066, 16'd771, 16'd54683, 16'd687, 16'd51169, 16'd58755}; // indx = 691
    #10;
    addra = 32'd22144;
    dina = {96'd0, 16'd50329, 16'd26635, 16'd26382, 16'd52304, 16'd46639, 16'd14621, 16'd64908, 16'd61971, 16'd33350, 16'd21633}; // indx = 692
    #10;
    addra = 32'd22176;
    dina = {96'd0, 16'd57478, 16'd17352, 16'd30154, 16'd35868, 16'd35836, 16'd3877, 16'd14746, 16'd30668, 16'd10548, 16'd22089}; // indx = 693
    #10;
    addra = 32'd22208;
    dina = {96'd0, 16'd18556, 16'd39617, 16'd60857, 16'd10478, 16'd16026, 16'd25729, 16'd26273, 16'd43104, 16'd24201, 16'd43190}; // indx = 694
    #10;
    addra = 32'd22240;
    dina = {96'd0, 16'd29243, 16'd38389, 16'd43859, 16'd38405, 16'd3576, 16'd1575, 16'd25631, 16'd30401, 16'd45136, 16'd31268}; // indx = 695
    #10;
    addra = 32'd22272;
    dina = {96'd0, 16'd24559, 16'd27063, 16'd43906, 16'd10362, 16'd19743, 16'd58304, 16'd49493, 16'd2464, 16'd37878, 16'd9136}; // indx = 696
    #10;
    addra = 32'd22304;
    dina = {96'd0, 16'd14539, 16'd13191, 16'd46976, 16'd59050, 16'd23144, 16'd44612, 16'd46005, 16'd22113, 16'd58816, 16'd27329}; // indx = 697
    #10;
    addra = 32'd22336;
    dina = {96'd0, 16'd58988, 16'd3198, 16'd40359, 16'd45002, 16'd10975, 16'd51171, 16'd39235, 16'd17182, 16'd18811, 16'd30997}; // indx = 698
    #10;
    addra = 32'd22368;
    dina = {96'd0, 16'd20973, 16'd7032, 16'd45695, 16'd19890, 16'd12392, 16'd36297, 16'd42793, 16'd9852, 16'd34495, 16'd57330}; // indx = 699
    #10;
    addra = 32'd22400;
    dina = {96'd0, 16'd63843, 16'd45231, 16'd25537, 16'd44608, 16'd38800, 16'd7126, 16'd51984, 16'd17506, 16'd61404, 16'd23636}; // indx = 700
    #10;
    addra = 32'd22432;
    dina = {96'd0, 16'd18101, 16'd31624, 16'd17013, 16'd53861, 16'd8133, 16'd48579, 16'd27874, 16'd16506, 16'd52451, 16'd21224}; // indx = 701
    #10;
    addra = 32'd22464;
    dina = {96'd0, 16'd55317, 16'd11675, 16'd696, 16'd34696, 16'd12670, 16'd29443, 16'd60047, 16'd52714, 16'd63257, 16'd43542}; // indx = 702
    #10;
    addra = 32'd22496;
    dina = {96'd0, 16'd57908, 16'd36050, 16'd47792, 16'd51624, 16'd26936, 16'd12843, 16'd24001, 16'd43244, 16'd13832, 16'd2600}; // indx = 703
    #10;
    addra = 32'd22528;
    dina = {96'd0, 16'd54906, 16'd58384, 16'd21603, 16'd728, 16'd32079, 16'd60214, 16'd45316, 16'd30674, 16'd6644, 16'd65081}; // indx = 704
    #10;
    addra = 32'd22560;
    dina = {96'd0, 16'd8109, 16'd13875, 16'd25016, 16'd14679, 16'd28244, 16'd35954, 16'd55035, 16'd32500, 16'd57732, 16'd58790}; // indx = 705
    #10;
    addra = 32'd22592;
    dina = {96'd0, 16'd53110, 16'd21959, 16'd17579, 16'd18020, 16'd57295, 16'd30877, 16'd21378, 16'd47422, 16'd24012, 16'd56492}; // indx = 706
    #10;
    addra = 32'd22624;
    dina = {96'd0, 16'd2279, 16'd13446, 16'd54345, 16'd7224, 16'd41975, 16'd39427, 16'd35952, 16'd36424, 16'd22702, 16'd30419}; // indx = 707
    #10;
    addra = 32'd22656;
    dina = {96'd0, 16'd20774, 16'd7092, 16'd48641, 16'd46548, 16'd38111, 16'd51962, 16'd1435, 16'd33473, 16'd25471, 16'd52789}; // indx = 708
    #10;
    addra = 32'd22688;
    dina = {96'd0, 16'd28665, 16'd10241, 16'd9521, 16'd39678, 16'd19119, 16'd1260, 16'd39629, 16'd10378, 16'd14377, 16'd23888}; // indx = 709
    #10;
    addra = 32'd22720;
    dina = {96'd0, 16'd53108, 16'd52108, 16'd19486, 16'd47321, 16'd49906, 16'd14352, 16'd32290, 16'd13847, 16'd5491, 16'd43153}; // indx = 710
    #10;
    addra = 32'd22752;
    dina = {96'd0, 16'd39251, 16'd56388, 16'd59823, 16'd7740, 16'd35219, 16'd36315, 16'd12594, 16'd20999, 16'd27674, 16'd62341}; // indx = 711
    #10;
    addra = 32'd22784;
    dina = {96'd0, 16'd47860, 16'd12964, 16'd19981, 16'd57460, 16'd46376, 16'd21219, 16'd20098, 16'd26428, 16'd26232, 16'd60626}; // indx = 712
    #10;
    addra = 32'd22816;
    dina = {96'd0, 16'd57362, 16'd4792, 16'd11344, 16'd46827, 16'd40161, 16'd4322, 16'd23788, 16'd53664, 16'd57801, 16'd44658}; // indx = 713
    #10;
    addra = 32'd22848;
    dina = {96'd0, 16'd15807, 16'd4388, 16'd30048, 16'd34033, 16'd51084, 16'd53360, 16'd57571, 16'd46568, 16'd21063, 16'd11148}; // indx = 714
    #10;
    addra = 32'd22880;
    dina = {96'd0, 16'd33085, 16'd17519, 16'd41389, 16'd8036, 16'd31078, 16'd35384, 16'd18786, 16'd47756, 16'd63269, 16'd25025}; // indx = 715
    #10;
    addra = 32'd22912;
    dina = {96'd0, 16'd2840, 16'd46807, 16'd61953, 16'd45296, 16'd6435, 16'd37126, 16'd9001, 16'd59450, 16'd34006, 16'd34404}; // indx = 716
    #10;
    addra = 32'd22944;
    dina = {96'd0, 16'd4927, 16'd9655, 16'd25523, 16'd60123, 16'd13209, 16'd29513, 16'd31446, 16'd37571, 16'd8250, 16'd63310}; // indx = 717
    #10;
    addra = 32'd22976;
    dina = {96'd0, 16'd25826, 16'd25390, 16'd38846, 16'd14869, 16'd7409, 16'd8986, 16'd49750, 16'd5791, 16'd43516, 16'd32019}; // indx = 718
    #10;
    addra = 32'd23008;
    dina = {96'd0, 16'd37543, 16'd30578, 16'd25393, 16'd41093, 16'd17366, 16'd34074, 16'd40366, 16'd38409, 16'd54665, 16'd39319}; // indx = 719
    #10;
    addra = 32'd23040;
    dina = {96'd0, 16'd29738, 16'd31929, 16'd55300, 16'd64820, 16'd11955, 16'd57734, 16'd43819, 16'd18208, 16'd32306, 16'd9419}; // indx = 720
    #10;
    addra = 32'd23072;
    dina = {96'd0, 16'd31466, 16'd60384, 16'd17488, 16'd58668, 16'd65327, 16'd22586, 16'd2486, 16'd30882, 16'd43739, 16'd12164}; // indx = 721
    #10;
    addra = 32'd23104;
    dina = {96'd0, 16'd7961, 16'd36206, 16'd21885, 16'd64098, 16'd60781, 16'd44098, 16'd47804, 16'd26096, 16'd33397, 16'd55065}; // indx = 722
    #10;
    addra = 32'd23136;
    dina = {96'd0, 16'd42373, 16'd64270, 16'd324, 16'd40867, 16'd60055, 16'd345, 16'd48796, 16'd24200, 16'd10813, 16'd55732}; // indx = 723
    #10;
    addra = 32'd23168;
    dina = {96'd0, 16'd9017, 16'd32847, 16'd41559, 16'd16057, 16'd60112, 16'd50721, 16'd37218, 16'd55876, 16'd2939, 16'd22811}; // indx = 724
    #10;
    addra = 32'd23200;
    dina = {96'd0, 16'd14740, 16'd14348, 16'd40262, 16'd25969, 16'd44099, 16'd46168, 16'd401, 16'd10088, 16'd44275, 16'd25351}; // indx = 725
    #10;
    addra = 32'd23232;
    dina = {96'd0, 16'd13835, 16'd19126, 16'd44090, 16'd44722, 16'd20058, 16'd26001, 16'd36966, 16'd46482, 16'd45759, 16'd51371}; // indx = 726
    #10;
    addra = 32'd23264;
    dina = {96'd0, 16'd33327, 16'd28485, 16'd14971, 16'd63762, 16'd60357, 16'd38732, 16'd17818, 16'd44811, 16'd40204, 16'd11390}; // indx = 727
    #10;
    addra = 32'd23296;
    dina = {96'd0, 16'd48517, 16'd61005, 16'd1821, 16'd21709, 16'd14143, 16'd24836, 16'd37169, 16'd48312, 16'd34125, 16'd34089}; // indx = 728
    #10;
    addra = 32'd23328;
    dina = {96'd0, 16'd30357, 16'd24150, 16'd27426, 16'd65077, 16'd24325, 16'd28742, 16'd38218, 16'd44846, 16'd27520, 16'd42202}; // indx = 729
    #10;
    addra = 32'd23360;
    dina = {96'd0, 16'd59008, 16'd28646, 16'd26157, 16'd30885, 16'd51394, 16'd21758, 16'd8470, 16'd27647, 16'd23392, 16'd6066}; // indx = 730
    #10;
    addra = 32'd23392;
    dina = {96'd0, 16'd3084, 16'd4667, 16'd58683, 16'd17997, 16'd6623, 16'd51000, 16'd13000, 16'd46104, 16'd30165, 16'd32621}; // indx = 731
    #10;
    addra = 32'd23424;
    dina = {96'd0, 16'd14845, 16'd45221, 16'd54973, 16'd59083, 16'd25249, 16'd20451, 16'd13716, 16'd12643, 16'd51866, 16'd44480}; // indx = 732
    #10;
    addra = 32'd23456;
    dina = {96'd0, 16'd41198, 16'd6189, 16'd23811, 16'd35741, 16'd35813, 16'd20011, 16'd11967, 16'd45642, 16'd36986, 16'd53479}; // indx = 733
    #10;
    addra = 32'd23488;
    dina = {96'd0, 16'd8449, 16'd12529, 16'd47055, 16'd60110, 16'd10400, 16'd18645, 16'd17486, 16'd12292, 16'd21873, 16'd46651}; // indx = 734
    #10;
    addra = 32'd23520;
    dina = {96'd0, 16'd25867, 16'd38012, 16'd44134, 16'd2897, 16'd21720, 16'd21373, 16'd12158, 16'd2181, 16'd9443, 16'd27852}; // indx = 735
    #10;
    addra = 32'd23552;
    dina = {96'd0, 16'd33448, 16'd32758, 16'd29347, 16'd31337, 16'd53857, 16'd47437, 16'd3143, 16'd5376, 16'd45694, 16'd31727}; // indx = 736
    #10;
    addra = 32'd23584;
    dina = {96'd0, 16'd21316, 16'd41724, 16'd47038, 16'd1090, 16'd65375, 16'd51342, 16'd10941, 16'd834, 16'd10999, 16'd15957}; // indx = 737
    #10;
    addra = 32'd23616;
    dina = {96'd0, 16'd57809, 16'd41709, 16'd36780, 16'd56194, 16'd8356, 16'd15351, 16'd37561, 16'd43040, 16'd35581, 16'd13218}; // indx = 738
    #10;
    addra = 32'd23648;
    dina = {96'd0, 16'd35522, 16'd48344, 16'd65406, 16'd37888, 16'd37341, 16'd64996, 16'd17729, 16'd56218, 16'd659, 16'd13883}; // indx = 739
    #10;
    addra = 32'd23680;
    dina = {96'd0, 16'd23442, 16'd16386, 16'd14042, 16'd210, 16'd47195, 16'd49138, 16'd32295, 16'd31367, 16'd7141, 16'd15019}; // indx = 740
    #10;
    addra = 32'd23712;
    dina = {96'd0, 16'd37009, 16'd21696, 16'd15465, 16'd55744, 16'd4199, 16'd19779, 16'd62768, 16'd18429, 16'd35504, 16'd18825}; // indx = 741
    #10;
    addra = 32'd23744;
    dina = {96'd0, 16'd20510, 16'd17649, 16'd45512, 16'd44902, 16'd38345, 16'd60665, 16'd45799, 16'd32662, 16'd17874, 16'd60127}; // indx = 742
    #10;
    addra = 32'd23776;
    dina = {96'd0, 16'd25992, 16'd1225, 16'd55962, 16'd28978, 16'd18168, 16'd10169, 16'd45218, 16'd46917, 16'd19905, 16'd10841}; // indx = 743
    #10;
    addra = 32'd23808;
    dina = {96'd0, 16'd3601, 16'd37368, 16'd52825, 16'd4417, 16'd12309, 16'd33634, 16'd50303, 16'd3509, 16'd15992, 16'd40871}; // indx = 744
    #10;
    addra = 32'd23840;
    dina = {96'd0, 16'd52511, 16'd58841, 16'd32538, 16'd52900, 16'd60868, 16'd48401, 16'd35670, 16'd5757, 16'd9506, 16'd46702}; // indx = 745
    #10;
    addra = 32'd23872;
    dina = {96'd0, 16'd10042, 16'd63643, 16'd60234, 16'd19243, 16'd22910, 16'd9737, 16'd64459, 16'd47924, 16'd21899, 16'd19815}; // indx = 746
    #10;
    addra = 32'd23904;
    dina = {96'd0, 16'd9900, 16'd19683, 16'd47960, 16'd2600, 16'd31947, 16'd52826, 16'd6682, 16'd9288, 16'd45134, 16'd6847}; // indx = 747
    #10;
    addra = 32'd23936;
    dina = {96'd0, 16'd2915, 16'd5721, 16'd50916, 16'd10557, 16'd14548, 16'd44320, 16'd32291, 16'd57417, 16'd57341, 16'd55417}; // indx = 748
    #10;
    addra = 32'd23968;
    dina = {96'd0, 16'd58704, 16'd39665, 16'd25602, 16'd39121, 16'd43390, 16'd12083, 16'd61354, 16'd19296, 16'd31376, 16'd4701}; // indx = 749
    #10;
    addra = 32'd24000;
    dina = {96'd0, 16'd31786, 16'd10772, 16'd58062, 16'd9627, 16'd48319, 16'd36532, 16'd1638, 16'd60515, 16'd10645, 16'd25709}; // indx = 750
    #10;
    addra = 32'd24032;
    dina = {96'd0, 16'd19936, 16'd15291, 16'd14137, 16'd36642, 16'd58491, 16'd58868, 16'd25359, 16'd55662, 16'd40401, 16'd32773}; // indx = 751
    #10;
    addra = 32'd24064;
    dina = {96'd0, 16'd1755, 16'd17325, 16'd3626, 16'd18796, 16'd55352, 16'd54144, 16'd9379, 16'd49122, 16'd30367, 16'd29945}; // indx = 752
    #10;
    addra = 32'd24096;
    dina = {96'd0, 16'd43072, 16'd50016, 16'd15662, 16'd13482, 16'd10251, 16'd52612, 16'd9666, 16'd18039, 16'd35631, 16'd44570}; // indx = 753
    #10;
    addra = 32'd24128;
    dina = {96'd0, 16'd5978, 16'd64674, 16'd36814, 16'd15550, 16'd50687, 16'd6926, 16'd20674, 16'd28108, 16'd59024, 16'd57591}; // indx = 754
    #10;
    addra = 32'd24160;
    dina = {96'd0, 16'd63473, 16'd16144, 16'd16463, 16'd10217, 16'd18464, 16'd56608, 16'd59546, 16'd28776, 16'd25730, 16'd32209}; // indx = 755
    #10;
    addra = 32'd24192;
    dina = {96'd0, 16'd45482, 16'd63899, 16'd21087, 16'd64136, 16'd60350, 16'd20358, 16'd17898, 16'd45033, 16'd63947, 16'd8306}; // indx = 756
    #10;
    addra = 32'd24224;
    dina = {96'd0, 16'd8234, 16'd4342, 16'd25851, 16'd29485, 16'd52375, 16'd11876, 16'd17910, 16'd312, 16'd5588, 16'd60743}; // indx = 757
    #10;
    addra = 32'd24256;
    dina = {96'd0, 16'd3199, 16'd59874, 16'd42757, 16'd37206, 16'd5082, 16'd42918, 16'd41381, 16'd3107, 16'd45256, 16'd28814}; // indx = 758
    #10;
    addra = 32'd24288;
    dina = {96'd0, 16'd35816, 16'd10482, 16'd16144, 16'd27277, 16'd62745, 16'd34204, 16'd21162, 16'd56674, 16'd29477, 16'd39937}; // indx = 759
    #10;
    addra = 32'd24320;
    dina = {96'd0, 16'd5764, 16'd28564, 16'd16419, 16'd14636, 16'd50438, 16'd15270, 16'd29492, 16'd48830, 16'd52347, 16'd60669}; // indx = 760
    #10;
    addra = 32'd24352;
    dina = {96'd0, 16'd58149, 16'd16654, 16'd51400, 16'd59698, 16'd26715, 16'd4999, 16'd41788, 16'd26684, 16'd38977, 16'd31497}; // indx = 761
    #10;
    addra = 32'd24384;
    dina = {96'd0, 16'd17150, 16'd25529, 16'd41731, 16'd28983, 16'd13847, 16'd15544, 16'd6778, 16'd48050, 16'd51506, 16'd64215}; // indx = 762
    #10;
    addra = 32'd24416;
    dina = {96'd0, 16'd44540, 16'd44967, 16'd13597, 16'd58534, 16'd40897, 16'd12308, 16'd9948, 16'd44608, 16'd423, 16'd29386}; // indx = 763
    #10;
    addra = 32'd24448;
    dina = {96'd0, 16'd26826, 16'd53806, 16'd36208, 16'd36006, 16'd25389, 16'd46097, 16'd50508, 16'd56716, 16'd14711, 16'd58432}; // indx = 764
    #10;
    addra = 32'd24480;
    dina = {96'd0, 16'd2992, 16'd32768, 16'd31012, 16'd30156, 16'd54526, 16'd37240, 16'd30432, 16'd63848, 16'd56997, 16'd45181}; // indx = 765
    #10;
    addra = 32'd24512;
    dina = {96'd0, 16'd20864, 16'd53375, 16'd54011, 16'd27215, 16'd22910, 16'd14528, 16'd58703, 16'd9994, 16'd26436, 16'd22350}; // indx = 766
    #10;
    addra = 32'd24544;
    dina = {96'd0, 16'd56744, 16'd38158, 16'd19916, 16'd17118, 16'd1204, 16'd12121, 16'd59410, 16'd4249, 16'd8197, 16'd36376}; // indx = 767
    #10;
    addra = 32'd24576;
    dina = {96'd0, 16'd29960, 16'd10942, 16'd40010, 16'd364, 16'd59561, 16'd7622, 16'd9152, 16'd4460, 16'd16741, 16'd24449}; // indx = 768
    #10;
    addra = 32'd24608;
    dina = {96'd0, 16'd3399, 16'd36949, 16'd31880, 16'd34765, 16'd32395, 16'd11100, 16'd21524, 16'd53988, 16'd29174, 16'd11017}; // indx = 769
    #10;
    addra = 32'd24640;
    dina = {96'd0, 16'd50455, 16'd25745, 16'd37144, 16'd58756, 16'd14265, 16'd32432, 16'd31545, 16'd45144, 16'd61784, 16'd2482}; // indx = 770
    #10;
    addra = 32'd24672;
    dina = {96'd0, 16'd54613, 16'd475, 16'd55592, 16'd18684, 16'd4399, 16'd13619, 16'd21367, 16'd19764, 16'd38120, 16'd9029}; // indx = 771
    #10;
    addra = 32'd24704;
    dina = {96'd0, 16'd5535, 16'd4617, 16'd33296, 16'd60321, 16'd31034, 16'd55461, 16'd51946, 16'd24014, 16'd17866, 16'd3850}; // indx = 772
    #10;
    addra = 32'd24736;
    dina = {96'd0, 16'd47629, 16'd32108, 16'd2531, 16'd21085, 16'd29030, 16'd21941, 16'd61775, 16'd19494, 16'd58261, 16'd15405}; // indx = 773
    #10;
    addra = 32'd24768;
    dina = {96'd0, 16'd12885, 16'd49691, 16'd63188, 16'd30527, 16'd46100, 16'd55449, 16'd42545, 16'd52156, 16'd11759, 16'd64104}; // indx = 774
    #10;
    addra = 32'd24800;
    dina = {96'd0, 16'd33353, 16'd26604, 16'd8033, 16'd59323, 16'd25868, 16'd49004, 16'd26625, 16'd39970, 16'd19291, 16'd46845}; // indx = 775
    #10;
    addra = 32'd24832;
    dina = {96'd0, 16'd1712, 16'd59446, 16'd35906, 16'd13567, 16'd776, 16'd53894, 16'd33876, 16'd5564, 16'd61227, 16'd55504}; // indx = 776
    #10;
    addra = 32'd24864;
    dina = {96'd0, 16'd28994, 16'd21402, 16'd10802, 16'd56834, 16'd56252, 16'd7076, 16'd30298, 16'd5661, 16'd63640, 16'd42544}; // indx = 777
    #10;
    addra = 32'd24896;
    dina = {96'd0, 16'd40506, 16'd4665, 16'd45669, 16'd34366, 16'd33917, 16'd6292, 16'd42972, 16'd37763, 16'd50482, 16'd26132}; // indx = 778
    #10;
    addra = 32'd24928;
    dina = {96'd0, 16'd8064, 16'd50487, 16'd47305, 16'd34440, 16'd58011, 16'd34070, 16'd58865, 16'd49342, 16'd60232, 16'd724}; // indx = 779
    #10;
    addra = 32'd24960;
    dina = {96'd0, 16'd24342, 16'd46758, 16'd61957, 16'd37094, 16'd59531, 16'd31988, 16'd25504, 16'd1073, 16'd37911, 16'd4847}; // indx = 780
    #10;
    addra = 32'd24992;
    dina = {96'd0, 16'd22413, 16'd11548, 16'd62363, 16'd65322, 16'd63625, 16'd12219, 16'd9878, 16'd55576, 16'd20880, 16'd1225}; // indx = 781
    #10;
    addra = 32'd25024;
    dina = {96'd0, 16'd37544, 16'd1961, 16'd42005, 16'd55428, 16'd41000, 16'd43380, 16'd25926, 16'd30621, 16'd7701, 16'd14978}; // indx = 782
    #10;
    addra = 32'd25056;
    dina = {96'd0, 16'd44623, 16'd31656, 16'd10772, 16'd11176, 16'd5237, 16'd61224, 16'd52486, 16'd60405, 16'd54233, 16'd21696}; // indx = 783
    #10;
    addra = 32'd25088;
    dina = {96'd0, 16'd5612, 16'd34786, 16'd13619, 16'd44289, 16'd29969, 16'd30367, 16'd48275, 16'd3977, 16'd9466, 16'd35657}; // indx = 784
    #10;
    addra = 32'd25120;
    dina = {96'd0, 16'd54840, 16'd6244, 16'd8055, 16'd42541, 16'd30268, 16'd8284, 16'd22358, 16'd41522, 16'd42852, 16'd43124}; // indx = 785
    #10;
    addra = 32'd25152;
    dina = {96'd0, 16'd58185, 16'd30969, 16'd58628, 16'd53712, 16'd47292, 16'd41881, 16'd36926, 16'd19849, 16'd35416, 16'd22265}; // indx = 786
    #10;
    addra = 32'd25184;
    dina = {96'd0, 16'd13390, 16'd22849, 16'd30886, 16'd14931, 16'd54600, 16'd1304, 16'd21908, 16'd51988, 16'd64485, 16'd37849}; // indx = 787
    #10;
    addra = 32'd25216;
    dina = {96'd0, 16'd64917, 16'd47523, 16'd60392, 16'd7214, 16'd38663, 16'd50579, 16'd24137, 16'd30069, 16'd10750, 16'd1922}; // indx = 788
    #10;
    addra = 32'd25248;
    dina = {96'd0, 16'd33303, 16'd2329, 16'd33631, 16'd11931, 16'd39947, 16'd18111, 16'd7049, 16'd55322, 16'd55062, 16'd10433}; // indx = 789
    #10;
    addra = 32'd25280;
    dina = {96'd0, 16'd6518, 16'd52739, 16'd46325, 16'd4384, 16'd2393, 16'd7443, 16'd41255, 16'd41807, 16'd9129, 16'd9710}; // indx = 790
    #10;
    addra = 32'd25312;
    dina = {96'd0, 16'd30889, 16'd14837, 16'd19788, 16'd41215, 16'd37417, 16'd63675, 16'd1572, 16'd59909, 16'd1872, 16'd45051}; // indx = 791
    #10;
    addra = 32'd25344;
    dina = {96'd0, 16'd18107, 16'd54917, 16'd3056, 16'd3565, 16'd54342, 16'd47535, 16'd15662, 16'd48278, 16'd49914, 16'd18731}; // indx = 792
    #10;
    addra = 32'd25376;
    dina = {96'd0, 16'd10231, 16'd11191, 16'd63451, 16'd36219, 16'd28235, 16'd6583, 16'd13190, 16'd32601, 16'd61285, 16'd614}; // indx = 793
    #10;
    addra = 32'd25408;
    dina = {96'd0, 16'd64658, 16'd12715, 16'd39329, 16'd29779, 16'd52861, 16'd21850, 16'd8736, 16'd56762, 16'd3280, 16'd42129}; // indx = 794
    #10;
    addra = 32'd25440;
    dina = {96'd0, 16'd14593, 16'd49638, 16'd60480, 16'd26238, 16'd4488, 16'd10863, 16'd55705, 16'd58982, 16'd50721, 16'd45497}; // indx = 795
    #10;
    addra = 32'd25472;
    dina = {96'd0, 16'd10313, 16'd49406, 16'd45776, 16'd17447, 16'd62148, 16'd11807, 16'd3455, 16'd21194, 16'd42921, 16'd55645}; // indx = 796
    #10;
    addra = 32'd25504;
    dina = {96'd0, 16'd56037, 16'd48481, 16'd47160, 16'd2247, 16'd64432, 16'd19220, 16'd51231, 16'd10548, 16'd50023, 16'd16387}; // indx = 797
    #10;
    addra = 32'd25536;
    dina = {96'd0, 16'd3112, 16'd38058, 16'd5222, 16'd22759, 16'd44136, 16'd63202, 16'd24674, 16'd30889, 16'd35718, 16'd27526}; // indx = 798
    #10;
    addra = 32'd25568;
    dina = {96'd0, 16'd64550, 16'd7599, 16'd19682, 16'd3443, 16'd42167, 16'd41910, 16'd40551, 16'd839, 16'd45561, 16'd35701}; // indx = 799
    #10;
    addra = 32'd25600;
    dina = {96'd0, 16'd12578, 16'd42822, 16'd50575, 16'd30089, 16'd34138, 16'd36619, 16'd60267, 16'd59498, 16'd4172, 16'd2709}; // indx = 800
    #10;
    addra = 32'd25632;
    dina = {96'd0, 16'd15023, 16'd52032, 16'd24588, 16'd20110, 16'd11936, 16'd34890, 16'd62800, 16'd50874, 16'd22909, 16'd21875}; // indx = 801
    #10;
    addra = 32'd25664;
    dina = {96'd0, 16'd6017, 16'd24135, 16'd22417, 16'd57366, 16'd59704, 16'd10062, 16'd61144, 16'd26219, 16'd1684, 16'd46871}; // indx = 802
    #10;
    addra = 32'd25696;
    dina = {96'd0, 16'd42482, 16'd47104, 16'd50475, 16'd35784, 16'd14985, 16'd7586, 16'd25837, 16'd9964, 16'd63636, 16'd59067}; // indx = 803
    #10;
    addra = 32'd25728;
    dina = {96'd0, 16'd27283, 16'd5868, 16'd40491, 16'd23242, 16'd17823, 16'd19864, 16'd41856, 16'd22147, 16'd29819, 16'd3575}; // indx = 804
    #10;
    addra = 32'd25760;
    dina = {96'd0, 16'd28543, 16'd29625, 16'd26385, 16'd50174, 16'd15949, 16'd44701, 16'd37917, 16'd7807, 16'd11750, 16'd7729}; // indx = 805
    #10;
    addra = 32'd25792;
    dina = {96'd0, 16'd15519, 16'd61294, 16'd48939, 16'd43596, 16'd41519, 16'd8755, 16'd48831, 16'd53893, 16'd44972, 16'd1966}; // indx = 806
    #10;
    addra = 32'd25824;
    dina = {96'd0, 16'd57966, 16'd44515, 16'd22810, 16'd50189, 16'd15793, 16'd28598, 16'd46444, 16'd33803, 16'd17148, 16'd42254}; // indx = 807
    #10;
    addra = 32'd25856;
    dina = {96'd0, 16'd29659, 16'd60505, 16'd55913, 16'd11119, 16'd44000, 16'd39177, 16'd31592, 16'd55657, 16'd44447, 16'd9704}; // indx = 808
    #10;
    addra = 32'd25888;
    dina = {96'd0, 16'd37529, 16'd49640, 16'd43968, 16'd13491, 16'd4505, 16'd48138, 16'd17839, 16'd49744, 16'd33717, 16'd54470}; // indx = 809
    #10;
    addra = 32'd25920;
    dina = {96'd0, 16'd50766, 16'd37192, 16'd36815, 16'd21021, 16'd19787, 16'd8762, 16'd10800, 16'd5814, 16'd310, 16'd11331}; // indx = 810
    #10;
    addra = 32'd25952;
    dina = {96'd0, 16'd58282, 16'd57602, 16'd38076, 16'd62448, 16'd7812, 16'd48561, 16'd21086, 16'd31354, 16'd18590, 16'd39969}; // indx = 811
    #10;
    addra = 32'd25984;
    dina = {96'd0, 16'd5568, 16'd15046, 16'd47835, 16'd35427, 16'd53119, 16'd50994, 16'd5847, 16'd14889, 16'd33030, 16'd2049}; // indx = 812
    #10;
    addra = 32'd26016;
    dina = {96'd0, 16'd19083, 16'd58584, 16'd4063, 16'd34785, 16'd11928, 16'd44224, 16'd58619, 16'd822, 16'd48047, 16'd34623}; // indx = 813
    #10;
    addra = 32'd26048;
    dina = {96'd0, 16'd47972, 16'd63370, 16'd35796, 16'd59050, 16'd46658, 16'd51656, 16'd49145, 16'd8833, 16'd3513, 16'd11604}; // indx = 814
    #10;
    addra = 32'd26080;
    dina = {96'd0, 16'd21713, 16'd43983, 16'd54178, 16'd18718, 16'd62688, 16'd11644, 16'd13660, 16'd32004, 16'd38382, 16'd20007}; // indx = 815
    #10;
    addra = 32'd26112;
    dina = {96'd0, 16'd38876, 16'd65199, 16'd23054, 16'd3216, 16'd57241, 16'd49871, 16'd15555, 16'd25204, 16'd57944, 16'd56176}; // indx = 816
    #10;
    addra = 32'd26144;
    dina = {96'd0, 16'd31366, 16'd20030, 16'd31815, 16'd10458, 16'd18088, 16'd28709, 16'd49391, 16'd2944, 16'd50538, 16'd19688}; // indx = 817
    #10;
    addra = 32'd26176;
    dina = {96'd0, 16'd59933, 16'd43567, 16'd41102, 16'd5779, 16'd50763, 16'd4994, 16'd49245, 16'd39547, 16'd113, 16'd60601}; // indx = 818
    #10;
    addra = 32'd26208;
    dina = {96'd0, 16'd26651, 16'd2721, 16'd22729, 16'd53674, 16'd16042, 16'd48646, 16'd29518, 16'd14602, 16'd38209, 16'd24348}; // indx = 819
    #10;
    addra = 32'd26240;
    dina = {96'd0, 16'd17391, 16'd47600, 16'd20590, 16'd31942, 16'd42739, 16'd19298, 16'd5163, 16'd8211, 16'd4299, 16'd39334}; // indx = 820
    #10;
    addra = 32'd26272;
    dina = {96'd0, 16'd28109, 16'd18198, 16'd41350, 16'd28142, 16'd16275, 16'd30076, 16'd33609, 16'd16749, 16'd9787, 16'd21904}; // indx = 821
    #10;
    addra = 32'd26304;
    dina = {96'd0, 16'd2179, 16'd51038, 16'd62377, 16'd49948, 16'd376, 16'd10957, 16'd49675, 16'd24777, 16'd64344, 16'd20443}; // indx = 822
    #10;
    addra = 32'd26336;
    dina = {96'd0, 16'd56355, 16'd44647, 16'd30207, 16'd11446, 16'd64986, 16'd7370, 16'd29629, 16'd57985, 16'd2795, 16'd57769}; // indx = 823
    #10;
    addra = 32'd26368;
    dina = {96'd0, 16'd15609, 16'd31882, 16'd64576, 16'd24842, 16'd23186, 16'd48020, 16'd2608, 16'd13678, 16'd26645, 16'd62396}; // indx = 824
    #10;
    addra = 32'd26400;
    dina = {96'd0, 16'd26074, 16'd8384, 16'd17627, 16'd50362, 16'd40279, 16'd48525, 16'd5758, 16'd17475, 16'd50724, 16'd34278}; // indx = 825
    #10;
    addra = 32'd26432;
    dina = {96'd0, 16'd60802, 16'd24045, 16'd33452, 16'd52650, 16'd32353, 16'd46559, 16'd54728, 16'd38518, 16'd21978, 16'd13599}; // indx = 826
    #10;
    addra = 32'd26464;
    dina = {96'd0, 16'd4621, 16'd19714, 16'd44010, 16'd44953, 16'd34562, 16'd7156, 16'd22040, 16'd36732, 16'd10938, 16'd47115}; // indx = 827
    #10;
    addra = 32'd26496;
    dina = {96'd0, 16'd35487, 16'd56212, 16'd9043, 16'd35492, 16'd53773, 16'd54672, 16'd49378, 16'd22590, 16'd18885, 16'd15487}; // indx = 828
    #10;
    addra = 32'd26528;
    dina = {96'd0, 16'd38395, 16'd9583, 16'd38391, 16'd63023, 16'd9774, 16'd62571, 16'd37410, 16'd9797, 16'd1647, 16'd44681}; // indx = 829
    #10;
    addra = 32'd26560;
    dina = {96'd0, 16'd23622, 16'd42187, 16'd3568, 16'd36565, 16'd19395, 16'd21804, 16'd48032, 16'd28912, 16'd16387, 16'd23491}; // indx = 830
    #10;
    addra = 32'd26592;
    dina = {96'd0, 16'd10679, 16'd24665, 16'd35454, 16'd19181, 16'd61451, 16'd57969, 16'd15803, 16'd27493, 16'd40643, 16'd28436}; // indx = 831
    #10;
    addra = 32'd26624;
    dina = {96'd0, 16'd3508, 16'd31698, 16'd37799, 16'd12159, 16'd22537, 16'd31803, 16'd36626, 16'd51424, 16'd36675, 16'd8132}; // indx = 832
    #10;
    addra = 32'd26656;
    dina = {96'd0, 16'd3364, 16'd14542, 16'd60014, 16'd10106, 16'd52277, 16'd23759, 16'd16229, 16'd41194, 16'd26704, 16'd48575}; // indx = 833
    #10;
    addra = 32'd26688;
    dina = {96'd0, 16'd54852, 16'd17750, 16'd53868, 16'd12102, 16'd38690, 16'd45414, 16'd7849, 16'd36963, 16'd61185, 16'd34092}; // indx = 834
    #10;
    addra = 32'd26720;
    dina = {96'd0, 16'd51856, 16'd37570, 16'd22757, 16'd33742, 16'd34625, 16'd58771, 16'd12823, 16'd23049, 16'd21878, 16'd16877}; // indx = 835
    #10;
    addra = 32'd26752;
    dina = {96'd0, 16'd32187, 16'd36481, 16'd12931, 16'd59895, 16'd11711, 16'd16187, 16'd45628, 16'd34821, 16'd12950, 16'd38566}; // indx = 836
    #10;
    addra = 32'd26784;
    dina = {96'd0, 16'd32785, 16'd27365, 16'd49876, 16'd48123, 16'd58726, 16'd54756, 16'd16944, 16'd2633, 16'd58817, 16'd13082}; // indx = 837
    #10;
    addra = 32'd26816;
    dina = {96'd0, 16'd59681, 16'd22757, 16'd39639, 16'd62546, 16'd24391, 16'd63780, 16'd8708, 16'd57950, 16'd57266, 16'd20058}; // indx = 838
    #10;
    addra = 32'd26848;
    dina = {96'd0, 16'd64984, 16'd15105, 16'd56770, 16'd33316, 16'd38025, 16'd6221, 16'd13475, 16'd60237, 16'd39750, 16'd6043}; // indx = 839
    #10;
    addra = 32'd26880;
    dina = {96'd0, 16'd4662, 16'd19670, 16'd19184, 16'd26395, 16'd33073, 16'd20144, 16'd16870, 16'd21151, 16'd44597, 16'd9697}; // indx = 840
    #10;
    addra = 32'd26912;
    dina = {96'd0, 16'd30392, 16'd55943, 16'd24636, 16'd7583, 16'd48235, 16'd31765, 16'd51065, 16'd29102, 16'd21530, 16'd48018}; // indx = 841
    #10;
    addra = 32'd26944;
    dina = {96'd0, 16'd37901, 16'd16224, 16'd56980, 16'd28577, 16'd2185, 16'd59883, 16'd34751, 16'd54580, 16'd63636, 16'd50287}; // indx = 842
    #10;
    addra = 32'd26976;
    dina = {96'd0, 16'd22834, 16'd12790, 16'd9689, 16'd17188, 16'd42055, 16'd27892, 16'd61195, 16'd54080, 16'd23770, 16'd50922}; // indx = 843
    #10;
    addra = 32'd27008;
    dina = {96'd0, 16'd21713, 16'd62793, 16'd547, 16'd62930, 16'd37611, 16'd42243, 16'd17959, 16'd58565, 16'd17183, 16'd33221}; // indx = 844
    #10;
    addra = 32'd27040;
    dina = {96'd0, 16'd31600, 16'd48975, 16'd27942, 16'd20196, 16'd58251, 16'd34325, 16'd27292, 16'd31634, 16'd47967, 16'd57567}; // indx = 845
    #10;
    addra = 32'd27072;
    dina = {96'd0, 16'd39622, 16'd44618, 16'd24349, 16'd64363, 16'd57476, 16'd2924, 16'd12674, 16'd55986, 16'd45542, 16'd19968}; // indx = 846
    #10;
    addra = 32'd27104;
    dina = {96'd0, 16'd2140, 16'd48775, 16'd137, 16'd33952, 16'd60218, 16'd25912, 16'd1046, 16'd3449, 16'd24747, 16'd10025}; // indx = 847
    #10;
    addra = 32'd27136;
    dina = {96'd0, 16'd43623, 16'd43595, 16'd15915, 16'd3485, 16'd64725, 16'd43675, 16'd2056, 16'd49383, 16'd31911, 16'd38544}; // indx = 848
    #10;
    addra = 32'd27168;
    dina = {96'd0, 16'd60287, 16'd22976, 16'd61240, 16'd24422, 16'd39836, 16'd55114, 16'd1941, 16'd4290, 16'd13925, 16'd54640}; // indx = 849
    #10;
    addra = 32'd27200;
    dina = {96'd0, 16'd58754, 16'd41649, 16'd61125, 16'd43142, 16'd45832, 16'd10341, 16'd64997, 16'd41849, 16'd21130, 16'd44044}; // indx = 850
    #10;
    addra = 32'd27232;
    dina = {96'd0, 16'd31381, 16'd52537, 16'd25085, 16'd57259, 16'd14821, 16'd43335, 16'd29780, 16'd1595, 16'd7937, 16'd39322}; // indx = 851
    #10;
    addra = 32'd27264;
    dina = {96'd0, 16'd53663, 16'd29882, 16'd25223, 16'd18695, 16'd47715, 16'd21668, 16'd33223, 16'd39783, 16'd52457, 16'd26263}; // indx = 852
    #10;
    addra = 32'd27296;
    dina = {96'd0, 16'd17693, 16'd8173, 16'd23527, 16'd61538, 16'd34321, 16'd23970, 16'd17257, 16'd32838, 16'd48528, 16'd27555}; // indx = 853
    #10;
    addra = 32'd27328;
    dina = {96'd0, 16'd53103, 16'd53362, 16'd7301, 16'd7245, 16'd28977, 16'd30589, 16'd9669, 16'd29788, 16'd16809, 16'd50582}; // indx = 854
    #10;
    addra = 32'd27360;
    dina = {96'd0, 16'd35104, 16'd31616, 16'd1894, 16'd37344, 16'd42063, 16'd64985, 16'd56431, 16'd21603, 16'd11871, 16'd8671}; // indx = 855
    #10;
    addra = 32'd27392;
    dina = {96'd0, 16'd54752, 16'd37476, 16'd47460, 16'd38106, 16'd26593, 16'd3787, 16'd21205, 16'd19080, 16'd14206, 16'd63602}; // indx = 856
    #10;
    addra = 32'd27424;
    dina = {96'd0, 16'd54354, 16'd37353, 16'd49019, 16'd39495, 16'd31870, 16'd11091, 16'd10091, 16'd14449, 16'd52542, 16'd40139}; // indx = 857
    #10;
    addra = 32'd27456;
    dina = {96'd0, 16'd12945, 16'd48330, 16'd8402, 16'd14079, 16'd37023, 16'd10537, 16'd10061, 16'd19144, 16'd43077, 16'd27652}; // indx = 858
    #10;
    addra = 32'd27488;
    dina = {96'd0, 16'd52161, 16'd44746, 16'd59442, 16'd2336, 16'd18276, 16'd25023, 16'd14316, 16'd64964, 16'd32279, 16'd40913}; // indx = 859
    #10;
    addra = 32'd27520;
    dina = {96'd0, 16'd8213, 16'd13027, 16'd44600, 16'd54481, 16'd43879, 16'd15049, 16'd48398, 16'd11124, 16'd35406, 16'd37265}; // indx = 860
    #10;
    addra = 32'd27552;
    dina = {96'd0, 16'd39316, 16'd30931, 16'd21619, 16'd18134, 16'd14456, 16'd16805, 16'd28897, 16'd28180, 16'd1431, 16'd61053}; // indx = 861
    #10;
    addra = 32'd27584;
    dina = {96'd0, 16'd25790, 16'd15313, 16'd4097, 16'd51478, 16'd22137, 16'd38768, 16'd33353, 16'd30636, 16'd12657, 16'd26222}; // indx = 862
    #10;
    addra = 32'd27616;
    dina = {96'd0, 16'd41188, 16'd14863, 16'd64659, 16'd13938, 16'd52792, 16'd48386, 16'd55792, 16'd2925, 16'd59015, 16'd35004}; // indx = 863
    #10;
    addra = 32'd27648;
    dina = {96'd0, 16'd63652, 16'd8251, 16'd26866, 16'd8597, 16'd42042, 16'd5238, 16'd56813, 16'd2956, 16'd38046, 16'd45996}; // indx = 864
    #10;
    addra = 32'd27680;
    dina = {96'd0, 16'd50961, 16'd21481, 16'd5188, 16'd15243, 16'd59080, 16'd49707, 16'd59510, 16'd17702, 16'd20891, 16'd65028}; // indx = 865
    #10;
    addra = 32'd27712;
    dina = {96'd0, 16'd41259, 16'd22950, 16'd28155, 16'd53318, 16'd15998, 16'd53138, 16'd29521, 16'd42704, 16'd2784, 16'd46615}; // indx = 866
    #10;
    addra = 32'd27744;
    dina = {96'd0, 16'd54267, 16'd38804, 16'd3533, 16'd40882, 16'd32646, 16'd22515, 16'd11391, 16'd50424, 16'd34314, 16'd5756}; // indx = 867
    #10;
    addra = 32'd27776;
    dina = {96'd0, 16'd11171, 16'd48577, 16'd2412, 16'd55414, 16'd58946, 16'd49303, 16'd10885, 16'd2867, 16'd47421, 16'd40678}; // indx = 868
    #10;
    addra = 32'd27808;
    dina = {96'd0, 16'd507, 16'd16128, 16'd49120, 16'd21910, 16'd10389, 16'd60917, 16'd55232, 16'd33589, 16'd27287, 16'd40530}; // indx = 869
    #10;
    addra = 32'd27840;
    dina = {96'd0, 16'd17165, 16'd4772, 16'd21939, 16'd19101, 16'd40917, 16'd18722, 16'd7871, 16'd17328, 16'd43527, 16'd1892}; // indx = 870
    #10;
    addra = 32'd27872;
    dina = {96'd0, 16'd1978, 16'd45829, 16'd27249, 16'd45895, 16'd34431, 16'd31558, 16'd3448, 16'd61870, 16'd24212, 16'd57310}; // indx = 871
    #10;
    addra = 32'd27904;
    dina = {96'd0, 16'd1197, 16'd9137, 16'd27282, 16'd63525, 16'd49078, 16'd31657, 16'd6796, 16'd44729, 16'd48390, 16'd37473}; // indx = 872
    #10;
    addra = 32'd27936;
    dina = {96'd0, 16'd54736, 16'd12702, 16'd3275, 16'd44352, 16'd47198, 16'd6494, 16'd53391, 16'd1428, 16'd38056, 16'd2287}; // indx = 873
    #10;
    addra = 32'd27968;
    dina = {96'd0, 16'd46009, 16'd44004, 16'd23148, 16'd35333, 16'd32504, 16'd18344, 16'd9815, 16'd12033, 16'd30833, 16'd44225}; // indx = 874
    #10;
    addra = 32'd28000;
    dina = {96'd0, 16'd17819, 16'd36174, 16'd17300, 16'd11103, 16'd60246, 16'd6169, 16'd42317, 16'd48148, 16'd26821, 16'd9908}; // indx = 875
    #10;
    addra = 32'd28032;
    dina = {96'd0, 16'd51662, 16'd24158, 16'd55942, 16'd30099, 16'd17239, 16'd40918, 16'd38048, 16'd28848, 16'd7421, 16'd11972}; // indx = 876
    #10;
    addra = 32'd28064;
    dina = {96'd0, 16'd27109, 16'd48491, 16'd10033, 16'd5754, 16'd48637, 16'd2907, 16'd15275, 16'd29661, 16'd41779, 16'd60381}; // indx = 877
    #10;
    addra = 32'd28096;
    dina = {96'd0, 16'd48975, 16'd50614, 16'd17976, 16'd56262, 16'd52281, 16'd17252, 16'd8475, 16'd8640, 16'd30176, 16'd30661}; // indx = 878
    #10;
    addra = 32'd28128;
    dina = {96'd0, 16'd36034, 16'd32307, 16'd63150, 16'd59142, 16'd4686, 16'd11470, 16'd58134, 16'd32601, 16'd37562, 16'd26368}; // indx = 879
    #10;
    addra = 32'd28160;
    dina = {96'd0, 16'd37201, 16'd38539, 16'd17164, 16'd59139, 16'd35760, 16'd53124, 16'd63998, 16'd56922, 16'd58382, 16'd26576}; // indx = 880
    #10;
    addra = 32'd28192;
    dina = {96'd0, 16'd36063, 16'd57175, 16'd25226, 16'd54513, 16'd39553, 16'd17687, 16'd48623, 16'd57072, 16'd33871, 16'd29584}; // indx = 881
    #10;
    addra = 32'd28224;
    dina = {96'd0, 16'd48183, 16'd47028, 16'd64705, 16'd53908, 16'd63851, 16'd17184, 16'd47690, 16'd38692, 16'd37610, 16'd22291}; // indx = 882
    #10;
    addra = 32'd28256;
    dina = {96'd0, 16'd20409, 16'd2436, 16'd26817, 16'd51379, 16'd50020, 16'd49987, 16'd5737, 16'd7230, 16'd16041, 16'd22617}; // indx = 883
    #10;
    addra = 32'd28288;
    dina = {96'd0, 16'd19236, 16'd53092, 16'd21443, 16'd49148, 16'd35676, 16'd61817, 16'd59948, 16'd32409, 16'd25358, 16'd47257}; // indx = 884
    #10;
    addra = 32'd28320;
    dina = {96'd0, 16'd52730, 16'd62879, 16'd54512, 16'd29915, 16'd10106, 16'd64601, 16'd45634, 16'd19525, 16'd63886, 16'd22553}; // indx = 885
    #10;
    addra = 32'd28352;
    dina = {96'd0, 16'd37033, 16'd11916, 16'd6272, 16'd27297, 16'd1056, 16'd39498, 16'd19299, 16'd22542, 16'd11213, 16'd19669}; // indx = 886
    #10;
    addra = 32'd28384;
    dina = {96'd0, 16'd47221, 16'd62998, 16'd44777, 16'd19444, 16'd14876, 16'd25889, 16'd51777, 16'd31880, 16'd53789, 16'd1272}; // indx = 887
    #10;
    addra = 32'd28416;
    dina = {96'd0, 16'd51324, 16'd38633, 16'd13613, 16'd17356, 16'd38955, 16'd6527, 16'd45809, 16'd22778, 16'd59553, 16'd1264}; // indx = 888
    #10;
    addra = 32'd28448;
    dina = {96'd0, 16'd63137, 16'd19072, 16'd9298, 16'd13173, 16'd17551, 16'd26476, 16'd58856, 16'd30168, 16'd14465, 16'd59841}; // indx = 889
    #10;
    addra = 32'd28480;
    dina = {96'd0, 16'd52353, 16'd44174, 16'd15753, 16'd58157, 16'd36695, 16'd57343, 16'd56804, 16'd44297, 16'd3762, 16'd63058}; // indx = 890
    #10;
    addra = 32'd28512;
    dina = {96'd0, 16'd64008, 16'd22372, 16'd3290, 16'd45365, 16'd4304, 16'd36013, 16'd24283, 16'd22887, 16'd30477, 16'd48522}; // indx = 891
    #10;
    addra = 32'd28544;
    dina = {96'd0, 16'd7600, 16'd15617, 16'd18215, 16'd31975, 16'd22694, 16'd49666, 16'd42911, 16'd43546, 16'd29438, 16'd64808}; // indx = 892
    #10;
    addra = 32'd28576;
    dina = {96'd0, 16'd48440, 16'd63232, 16'd60432, 16'd14240, 16'd10805, 16'd18939, 16'd16883, 16'd41063, 16'd43557, 16'd50896}; // indx = 893
    #10;
    addra = 32'd28608;
    dina = {96'd0, 16'd9113, 16'd33106, 16'd1657, 16'd2728, 16'd39211, 16'd29491, 16'd21807, 16'd43975, 16'd64515, 16'd1309}; // indx = 894
    #10;
    addra = 32'd28640;
    dina = {96'd0, 16'd56650, 16'd35811, 16'd32619, 16'd15172, 16'd44227, 16'd52499, 16'd48355, 16'd7653, 16'd43862, 16'd28668}; // indx = 895
    #10;
    addra = 32'd28672;
    dina = {96'd0, 16'd39239, 16'd7112, 16'd54583, 16'd57326, 16'd62284, 16'd6219, 16'd63426, 16'd13280, 16'd39712, 16'd19262}; // indx = 896
    #10;
    addra = 32'd28704;
    dina = {96'd0, 16'd40146, 16'd60689, 16'd53766, 16'd53533, 16'd27609, 16'd12334, 16'd16313, 16'd54077, 16'd40338, 16'd58671}; // indx = 897
    #10;
    addra = 32'd28736;
    dina = {96'd0, 16'd37205, 16'd42589, 16'd53386, 16'd25004, 16'd35878, 16'd45024, 16'd31859, 16'd25380, 16'd34061, 16'd53798}; // indx = 898
    #10;
    addra = 32'd28768;
    dina = {96'd0, 16'd64321, 16'd49595, 16'd43703, 16'd61260, 16'd54678, 16'd48157, 16'd29339, 16'd4907, 16'd62400, 16'd26278}; // indx = 899
    #10;
    addra = 32'd28800;
    dina = {96'd0, 16'd1277, 16'd4601, 16'd14328, 16'd33717, 16'd37873, 16'd22385, 16'd59276, 16'd31838, 16'd38813, 16'd22867}; // indx = 900
    #10;
    addra = 32'd28832;
    dina = {96'd0, 16'd13283, 16'd17601, 16'd25404, 16'd45397, 16'd23128, 16'd42039, 16'd22259, 16'd56116, 16'd39251, 16'd23608}; // indx = 901
    #10;
    addra = 32'd28864;
    dina = {96'd0, 16'd16606, 16'd33404, 16'd34963, 16'd49788, 16'd7190, 16'd55769, 16'd55999, 16'd16875, 16'd43382, 16'd7064}; // indx = 902
    #10;
    addra = 32'd28896;
    dina = {96'd0, 16'd44594, 16'd28163, 16'd63226, 16'd45781, 16'd30189, 16'd61030, 16'd26418, 16'd47646, 16'd59007, 16'd7281}; // indx = 903
    #10;
    addra = 32'd28928;
    dina = {96'd0, 16'd62673, 16'd32544, 16'd17870, 16'd61805, 16'd36025, 16'd16066, 16'd14107, 16'd51005, 16'd15803, 16'd10462}; // indx = 904
    #10;
    addra = 32'd28960;
    dina = {96'd0, 16'd62932, 16'd20634, 16'd25271, 16'd64653, 16'd24467, 16'd39705, 16'd4399, 16'd7849, 16'd14568, 16'd12118}; // indx = 905
    #10;
    addra = 32'd28992;
    dina = {96'd0, 16'd39323, 16'd47381, 16'd20531, 16'd2263, 16'd25916, 16'd21261, 16'd50141, 16'd6718, 16'd65461, 16'd29500}; // indx = 906
    #10;
    addra = 32'd29024;
    dina = {96'd0, 16'd7577, 16'd47469, 16'd5204, 16'd58095, 16'd56039, 16'd18036, 16'd12396, 16'd47092, 16'd21953, 16'd12649}; // indx = 907
    #10;
    addra = 32'd29056;
    dina = {96'd0, 16'd33100, 16'd6969, 16'd9738, 16'd34691, 16'd57267, 16'd62610, 16'd65182, 16'd41795, 16'd37458, 16'd64607}; // indx = 908
    #10;
    addra = 32'd29088;
    dina = {96'd0, 16'd14287, 16'd48108, 16'd41149, 16'd17231, 16'd51945, 16'd31999, 16'd55323, 16'd55618, 16'd52146, 16'd30847}; // indx = 909
    #10;
    addra = 32'd29120;
    dina = {96'd0, 16'd17225, 16'd46408, 16'd64081, 16'd12355, 16'd61718, 16'd49339, 16'd26331, 16'd10552, 16'd13316, 16'd9163}; // indx = 910
    #10;
    addra = 32'd29152;
    dina = {96'd0, 16'd26665, 16'd47874, 16'd59069, 16'd56304, 16'd37410, 16'd36626, 16'd63006, 16'd9633, 16'd23267, 16'd22390}; // indx = 911
    #10;
    addra = 32'd29184;
    dina = {96'd0, 16'd55438, 16'd22709, 16'd61748, 16'd28069, 16'd2338, 16'd18619, 16'd39708, 16'd7281, 16'd34054, 16'd50640}; // indx = 912
    #10;
    addra = 32'd29216;
    dina = {96'd0, 16'd30757, 16'd55635, 16'd31687, 16'd1072, 16'd25446, 16'd3613, 16'd40480, 16'd12522, 16'd30649, 16'd9226}; // indx = 913
    #10;
    addra = 32'd29248;
    dina = {96'd0, 16'd20163, 16'd47889, 16'd62447, 16'd4550, 16'd24574, 16'd10900, 16'd4735, 16'd54813, 16'd59905, 16'd25940}; // indx = 914
    #10;
    addra = 32'd29280;
    dina = {96'd0, 16'd9283, 16'd61717, 16'd10321, 16'd40343, 16'd42919, 16'd43370, 16'd50525, 16'd48565, 16'd34482, 16'd15859}; // indx = 915
    #10;
    addra = 32'd29312;
    dina = {96'd0, 16'd64712, 16'd19300, 16'd41152, 16'd28702, 16'd14758, 16'd41028, 16'd24780, 16'd4996, 16'd22290, 16'd64844}; // indx = 916
    #10;
    addra = 32'd29344;
    dina = {96'd0, 16'd43154, 16'd25302, 16'd45124, 16'd6803, 16'd6762, 16'd64913, 16'd15740, 16'd61238, 16'd56690, 16'd5488}; // indx = 917
    #10;
    addra = 32'd29376;
    dina = {96'd0, 16'd33797, 16'd37420, 16'd63943, 16'd58594, 16'd24799, 16'd44850, 16'd56743, 16'd2275, 16'd57386, 16'd37198}; // indx = 918
    #10;
    addra = 32'd29408;
    dina = {96'd0, 16'd83, 16'd3976, 16'd55504, 16'd19263, 16'd52634, 16'd16022, 16'd15914, 16'd5830, 16'd51593, 16'd18099}; // indx = 919
    #10;
    addra = 32'd29440;
    dina = {96'd0, 16'd14039, 16'd41839, 16'd35293, 16'd14911, 16'd5360, 16'd36151, 16'd32522, 16'd24439, 16'd52691, 16'd38582}; // indx = 920
    #10;
    addra = 32'd29472;
    dina = {96'd0, 16'd59032, 16'd17560, 16'd39718, 16'd35074, 16'd42603, 16'd62591, 16'd5841, 16'd34755, 16'd45050, 16'd61065}; // indx = 921
    #10;
    addra = 32'd29504;
    dina = {96'd0, 16'd43020, 16'd22265, 16'd21880, 16'd24060, 16'd10137, 16'd43353, 16'd55651, 16'd62589, 16'd1584, 16'd9635}; // indx = 922
    #10;
    addra = 32'd29536;
    dina = {96'd0, 16'd16991, 16'd42869, 16'd46913, 16'd17893, 16'd10104, 16'd36104, 16'd44090, 16'd44132, 16'd10899, 16'd3730}; // indx = 923
    #10;
    addra = 32'd29568;
    dina = {96'd0, 16'd39452, 16'd18117, 16'd30725, 16'd22031, 16'd61133, 16'd38821, 16'd20513, 16'd7932, 16'd60505, 16'd25734}; // indx = 924
    #10;
    addra = 32'd29600;
    dina = {96'd0, 16'd2717, 16'd45145, 16'd751, 16'd22937, 16'd19412, 16'd10616, 16'd38560, 16'd9990, 16'd54535, 16'd46380}; // indx = 925
    #10;
    addra = 32'd29632;
    dina = {96'd0, 16'd15020, 16'd57900, 16'd22112, 16'd61251, 16'd53593, 16'd45581, 16'd41730, 16'd27417, 16'd55535, 16'd59814}; // indx = 926
    #10;
    addra = 32'd29664;
    dina = {96'd0, 16'd22897, 16'd65050, 16'd6298, 16'd55161, 16'd62177, 16'd12901, 16'd55715, 16'd28676, 16'd32802, 16'd32904}; // indx = 927
    #10;
    addra = 32'd29696;
    dina = {96'd0, 16'd52884, 16'd22540, 16'd12324, 16'd1125, 16'd46919, 16'd3470, 16'd56822, 16'd37105, 16'd56614, 16'd4719}; // indx = 928
    #10;
    addra = 32'd29728;
    dina = {96'd0, 16'd26718, 16'd20922, 16'd34908, 16'd46104, 16'd32800, 16'd35854, 16'd29253, 16'd57739, 16'd50926, 16'd11472}; // indx = 929
    #10;
    addra = 32'd29760;
    dina = {96'd0, 16'd9098, 16'd38725, 16'd30961, 16'd1690, 16'd33307, 16'd23453, 16'd5420, 16'd39157, 16'd3588, 16'd43061}; // indx = 930
    #10;
    addra = 32'd29792;
    dina = {96'd0, 16'd38215, 16'd24474, 16'd34010, 16'd14871, 16'd43366, 16'd30856, 16'd22262, 16'd41830, 16'd55122, 16'd10622}; // indx = 931
    #10;
    addra = 32'd29824;
    dina = {96'd0, 16'd3047, 16'd8435, 16'd20481, 16'd30633, 16'd49332, 16'd31024, 16'd44063, 16'd5817, 16'd64991, 16'd47359}; // indx = 932
    #10;
    addra = 32'd29856;
    dina = {96'd0, 16'd50443, 16'd31766, 16'd38132, 16'd65416, 16'd28349, 16'd30449, 16'd24241, 16'd106, 16'd51518, 16'd14097}; // indx = 933
    #10;
    addra = 32'd29888;
    dina = {96'd0, 16'd61393, 16'd21056, 16'd35420, 16'd30986, 16'd38999, 16'd7121, 16'd64053, 16'd53424, 16'd32064, 16'd44943}; // indx = 934
    #10;
    addra = 32'd29920;
    dina = {96'd0, 16'd58977, 16'd8708, 16'd39443, 16'd3257, 16'd35678, 16'd45139, 16'd26009, 16'd31276, 16'd5789, 16'd58440}; // indx = 935
    #10;
    addra = 32'd29952;
    dina = {96'd0, 16'd10595, 16'd14517, 16'd2016, 16'd51338, 16'd58364, 16'd29296, 16'd54641, 16'd51547, 16'd1204, 16'd6491}; // indx = 936
    #10;
    addra = 32'd29984;
    dina = {96'd0, 16'd65293, 16'd60692, 16'd42169, 16'd33490, 16'd26415, 16'd58703, 16'd1888, 16'd57891, 16'd55417, 16'd61743}; // indx = 937
    #10;
    addra = 32'd30016;
    dina = {96'd0, 16'd49753, 16'd44298, 16'd12520, 16'd671, 16'd21821, 16'd57041, 16'd58977, 16'd47583, 16'd44293, 16'd31113}; // indx = 938
    #10;
    addra = 32'd30048;
    dina = {96'd0, 16'd64761, 16'd15515, 16'd22749, 16'd49057, 16'd32606, 16'd33393, 16'd5133, 16'd53863, 16'd3306, 16'd20309}; // indx = 939
    #10;
    addra = 32'd30080;
    dina = {96'd0, 16'd36167, 16'd31814, 16'd13063, 16'd47860, 16'd45005, 16'd4750, 16'd7557, 16'd18000, 16'd509, 16'd64411}; // indx = 940
    #10;
    addra = 32'd30112;
    dina = {96'd0, 16'd39086, 16'd5811, 16'd19957, 16'd52433, 16'd8628, 16'd8616, 16'd63689, 16'd54447, 16'd60828, 16'd39456}; // indx = 941
    #10;
    addra = 32'd30144;
    dina = {96'd0, 16'd3222, 16'd35632, 16'd43800, 16'd53444, 16'd59643, 16'd28894, 16'd40334, 16'd2466, 16'd18099, 16'd3502}; // indx = 942
    #10;
    addra = 32'd30176;
    dina = {96'd0, 16'd62797, 16'd38836, 16'd29889, 16'd45266, 16'd27505, 16'd50715, 16'd28459, 16'd28447, 16'd36380, 16'd43220}; // indx = 943
    #10;
    addra = 32'd30208;
    dina = {96'd0, 16'd59542, 16'd62361, 16'd40674, 16'd29182, 16'd9208, 16'd13542, 16'd3052, 16'd1263, 16'd23709, 16'd44073}; // indx = 944
    #10;
    addra = 32'd30240;
    dina = {96'd0, 16'd12550, 16'd45339, 16'd1396, 16'd9665, 16'd18073, 16'd5508, 16'd22085, 16'd23469, 16'd63566, 16'd41259}; // indx = 945
    #10;
    addra = 32'd30272;
    dina = {96'd0, 16'd39432, 16'd18211, 16'd41136, 16'd4235, 16'd55008, 16'd29685, 16'd45570, 16'd36785, 16'd6502, 16'd34736}; // indx = 946
    #10;
    addra = 32'd30304;
    dina = {96'd0, 16'd50471, 16'd55275, 16'd38201, 16'd17060, 16'd14499, 16'd41061, 16'd52107, 16'd50081, 16'd33425, 16'd59970}; // indx = 947
    #10;
    addra = 32'd30336;
    dina = {96'd0, 16'd43455, 16'd16337, 16'd27402, 16'd11526, 16'd30381, 16'd19099, 16'd9523, 16'd42413, 16'd8681, 16'd5554}; // indx = 948
    #10;
    addra = 32'd30368;
    dina = {96'd0, 16'd12714, 16'd47276, 16'd47978, 16'd31971, 16'd33544, 16'd7388, 16'd29594, 16'd51711, 16'd52691, 16'd34385}; // indx = 949
    #10;
    addra = 32'd30400;
    dina = {96'd0, 16'd19388, 16'd45913, 16'd11852, 16'd29796, 16'd13558, 16'd27123, 16'd6422, 16'd44466, 16'd44632, 16'd5176}; // indx = 950
    #10;
    addra = 32'd30432;
    dina = {96'd0, 16'd35002, 16'd17750, 16'd8077, 16'd3645, 16'd42096, 16'd23588, 16'd3045, 16'd3387, 16'd377, 16'd23546}; // indx = 951
    #10;
    addra = 32'd30464;
    dina = {96'd0, 16'd46523, 16'd1010, 16'd63675, 16'd32973, 16'd51654, 16'd50726, 16'd56156, 16'd64048, 16'd42307, 16'd44365}; // indx = 952
    #10;
    addra = 32'd30496;
    dina = {96'd0, 16'd5325, 16'd12737, 16'd2225, 16'd17363, 16'd37067, 16'd4014, 16'd38159, 16'd10187, 16'd48519, 16'd2313}; // indx = 953
    #10;
    addra = 32'd30528;
    dina = {96'd0, 16'd39026, 16'd27331, 16'd8445, 16'd31370, 16'd58705, 16'd61493, 16'd5320, 16'd18181, 16'd36338, 16'd21421}; // indx = 954
    #10;
    addra = 32'd30560;
    dina = {96'd0, 16'd9976, 16'd3433, 16'd15198, 16'd57321, 16'd29077, 16'd60282, 16'd41887, 16'd28977, 16'd60562, 16'd46019}; // indx = 955
    #10;
    addra = 32'd30592;
    dina = {96'd0, 16'd987, 16'd17872, 16'd9626, 16'd17046, 16'd6035, 16'd22047, 16'd45865, 16'd57301, 16'd59034, 16'd2425}; // indx = 956
    #10;
    addra = 32'd30624;
    dina = {96'd0, 16'd64179, 16'd22975, 16'd53681, 16'd14478, 16'd63833, 16'd6203, 16'd25704, 16'd62915, 16'd16200, 16'd38331}; // indx = 957
    #10;
    addra = 32'd30656;
    dina = {96'd0, 16'd35539, 16'd39957, 16'd38081, 16'd52504, 16'd25276, 16'd3713, 16'd42370, 16'd58175, 16'd19150, 16'd4035}; // indx = 958
    #10;
    addra = 32'd30688;
    dina = {96'd0, 16'd42698, 16'd28278, 16'd18405, 16'd50989, 16'd25246, 16'd40335, 16'd62352, 16'd43181, 16'd30844, 16'd6021}; // indx = 959
    #10;
    addra = 32'd30720;
    dina = {96'd0, 16'd21675, 16'd20236, 16'd53391, 16'd13839, 16'd27105, 16'd52644, 16'd8525, 16'd56037, 16'd35155, 16'd35520}; // indx = 960
    #10;
    addra = 32'd30752;
    dina = {96'd0, 16'd36389, 16'd29255, 16'd13615, 16'd31228, 16'd51443, 16'd49266, 16'd49473, 16'd53611, 16'd54621, 16'd28147}; // indx = 961
    #10;
    addra = 32'd30784;
    dina = {96'd0, 16'd45548, 16'd46291, 16'd51146, 16'd30809, 16'd7168, 16'd53935, 16'd52307, 16'd49975, 16'd21020, 16'd26954}; // indx = 962
    #10;
    addra = 32'd30816;
    dina = {96'd0, 16'd14222, 16'd24562, 16'd16902, 16'd40927, 16'd6624, 16'd47090, 16'd63286, 16'd19139, 16'd10411, 16'd6572}; // indx = 963
    #10;
    addra = 32'd30848;
    dina = {96'd0, 16'd24815, 16'd43421, 16'd12795, 16'd45877, 16'd9784, 16'd17511, 16'd43668, 16'd5769, 16'd34377, 16'd50656}; // indx = 964
    #10;
    addra = 32'd30880;
    dina = {96'd0, 16'd50469, 16'd4011, 16'd1789, 16'd54366, 16'd49672, 16'd52665, 16'd26997, 16'd59011, 16'd56337, 16'd62397}; // indx = 965
    #10;
    addra = 32'd30912;
    dina = {96'd0, 16'd14870, 16'd7589, 16'd54039, 16'd31961, 16'd3572, 16'd22488, 16'd19279, 16'd48970, 16'd27802, 16'd45991}; // indx = 966
    #10;
    addra = 32'd30944;
    dina = {96'd0, 16'd2210, 16'd13012, 16'd64305, 16'd29195, 16'd19539, 16'd9873, 16'd46429, 16'd48566, 16'd51527, 16'd16632}; // indx = 967
    #10;
    addra = 32'd30976;
    dina = {96'd0, 16'd64445, 16'd55095, 16'd37477, 16'd32678, 16'd3174, 16'd30310, 16'd34432, 16'd42460, 16'd10732, 16'd42911}; // indx = 968
    #10;
    addra = 32'd31008;
    dina = {96'd0, 16'd13552, 16'd7501, 16'd42704, 16'd56235, 16'd28614, 16'd58395, 16'd61682, 16'd46032, 16'd9072, 16'd44276}; // indx = 969
    #10;
    addra = 32'd31040;
    dina = {96'd0, 16'd48871, 16'd31106, 16'd30706, 16'd64383, 16'd29877, 16'd14729, 16'd5083, 16'd1389, 16'd36610, 16'd4135}; // indx = 970
    #10;
    addra = 32'd31072;
    dina = {96'd0, 16'd26288, 16'd41366, 16'd11436, 16'd50609, 16'd355, 16'd33902, 16'd18603, 16'd10, 16'd42331, 16'd65167}; // indx = 971
    #10;
    addra = 32'd31104;
    dina = {96'd0, 16'd9815, 16'd22956, 16'd20043, 16'd4983, 16'd18450, 16'd4705, 16'd5904, 16'd44630, 16'd2799, 16'd40489}; // indx = 972
    #10;
    addra = 32'd31136;
    dina = {96'd0, 16'd22948, 16'd26833, 16'd12399, 16'd21968, 16'd37965, 16'd34927, 16'd22611, 16'd21786, 16'd3802, 16'd11291}; // indx = 973
    #10;
    addra = 32'd31168;
    dina = {96'd0, 16'd43419, 16'd9410, 16'd59059, 16'd211, 16'd26941, 16'd6974, 16'd21764, 16'd46266, 16'd38255, 16'd48902}; // indx = 974
    #10;
    addra = 32'd31200;
    dina = {96'd0, 16'd8924, 16'd53652, 16'd50082, 16'd2218, 16'd28, 16'd6826, 16'd20208, 16'd64768, 16'd49114, 16'd8518}; // indx = 975
    #10;
    addra = 32'd31232;
    dina = {96'd0, 16'd2082, 16'd51578, 16'd54386, 16'd34292, 16'd3797, 16'd21015, 16'd4054, 16'd62332, 16'd43196, 16'd56315}; // indx = 976
    #10;
    addra = 32'd31264;
    dina = {96'd0, 16'd56832, 16'd9472, 16'd7574, 16'd32064, 16'd32988, 16'd41160, 16'd44884, 16'd59859, 16'd2499, 16'd48821}; // indx = 977
    #10;
    addra = 32'd31296;
    dina = {96'd0, 16'd20550, 16'd10520, 16'd9309, 16'd39768, 16'd41006, 16'd45599, 16'd50393, 16'd30853, 16'd29813, 16'd55720}; // indx = 978
    #10;
    addra = 32'd31328;
    dina = {96'd0, 16'd12702, 16'd30128, 16'd42158, 16'd62783, 16'd30387, 16'd34529, 16'd35989, 16'd28627, 16'd57232, 16'd29488}; // indx = 979
    #10;
    addra = 32'd31360;
    dina = {96'd0, 16'd56496, 16'd54907, 16'd56299, 16'd33891, 16'd40959, 16'd28572, 16'd38029, 16'd60568, 16'd17612, 16'd9742}; // indx = 980
    #10;
    addra = 32'd31392;
    dina = {96'd0, 16'd32445, 16'd56217, 16'd10347, 16'd4252, 16'd1836, 16'd14887, 16'd3245, 16'd33549, 16'd38293, 16'd63683}; // indx = 981
    #10;
    addra = 32'd31424;
    dina = {96'd0, 16'd31981, 16'd27735, 16'd36608, 16'd54176, 16'd64733, 16'd44892, 16'd21341, 16'd58903, 16'd63407, 16'd38401}; // indx = 982
    #10;
    addra = 32'd31456;
    dina = {96'd0, 16'd25871, 16'd392, 16'd62246, 16'd12173, 16'd60747, 16'd45825, 16'd46746, 16'd34632, 16'd12664, 16'd14539}; // indx = 983
    #10;
    addra = 32'd31488;
    dina = {96'd0, 16'd42444, 16'd2801, 16'd10398, 16'd28124, 16'd35457, 16'd64917, 16'd4713, 16'd65491, 16'd18019, 16'd58994}; // indx = 984
    #10;
    addra = 32'd31520;
    dina = {96'd0, 16'd17595, 16'd7944, 16'd58695, 16'd43675, 16'd19616, 16'd44721, 16'd41021, 16'd11582, 16'd21325, 16'd54433}; // indx = 985
    #10;
    addra = 32'd31552;
    dina = {96'd0, 16'd18292, 16'd17901, 16'd10049, 16'd55592, 16'd25733, 16'd2981, 16'd51723, 16'd8316, 16'd60019, 16'd11702}; // indx = 986
    #10;
    addra = 32'd31584;
    dina = {96'd0, 16'd10473, 16'd64307, 16'd9231, 16'd46851, 16'd32257, 16'd19727, 16'd63090, 16'd7633, 16'd15446, 16'd61926}; // indx = 987
    #10;
    addra = 32'd31616;
    dina = {96'd0, 16'd53108, 16'd19161, 16'd4539, 16'd52267, 16'd50364, 16'd39269, 16'd65256, 16'd22851, 16'd38937, 16'd19573}; // indx = 988
    #10;
    addra = 32'd31648;
    dina = {96'd0, 16'd42279, 16'd37861, 16'd60783, 16'd16213, 16'd64280, 16'd63057, 16'd35569, 16'd341, 16'd13807, 16'd34064}; // indx = 989
    #10;
    addra = 32'd31680;
    dina = {96'd0, 16'd52159, 16'd47851, 16'd59294, 16'd14633, 16'd16360, 16'd56312, 16'd6654, 16'd11058, 16'd32008, 16'd60363}; // indx = 990
    #10;
    addra = 32'd31712;
    dina = {96'd0, 16'd32570, 16'd60452, 16'd16862, 16'd50523, 16'd52845, 16'd62283, 16'd7561, 16'd53337, 16'd65374, 16'd22081}; // indx = 991
    #10;
    addra = 32'd31744;
    dina = {96'd0, 16'd8804, 16'd64959, 16'd58745, 16'd3880, 16'd44897, 16'd47557, 16'd2302, 16'd25757, 16'd62660, 16'd6371}; // indx = 992
    #10;
    addra = 32'd31776;
    dina = {96'd0, 16'd46535, 16'd34698, 16'd25413, 16'd8876, 16'd36639, 16'd12706, 16'd10155, 16'd3314, 16'd31862, 16'd50969}; // indx = 993
    #10;
    addra = 32'd31808;
    dina = {96'd0, 16'd47643, 16'd15379, 16'd34867, 16'd2599, 16'd37515, 16'd4838, 16'd32528, 16'd5194, 16'd13104, 16'd6537}; // indx = 994
    #10;
    addra = 32'd31840;
    dina = {96'd0, 16'd2361, 16'd10576, 16'd41012, 16'd60468, 16'd47074, 16'd44527, 16'd48702, 16'd35537, 16'd57579, 16'd65414}; // indx = 995
    #10;
    addra = 32'd31872;
    dina = {96'd0, 16'd45550, 16'd36868, 16'd64293, 16'd13046, 16'd37221, 16'd15385, 16'd16632, 16'd49211, 16'd46438, 16'd35332}; // indx = 996
    #10;
    addra = 32'd31904;
    dina = {96'd0, 16'd37377, 16'd14010, 16'd26909, 16'd46790, 16'd16219, 16'd46035, 16'd12523, 16'd12365, 16'd41812, 16'd51043}; // indx = 997
    #10;
    addra = 32'd31936;
    dina = {96'd0, 16'd13056, 16'd4160, 16'd44515, 16'd30601, 16'd14088, 16'd24700, 16'd5491, 16'd29476, 16'd26584, 16'd54787}; // indx = 998
    #10;
    addra = 32'd31968;
    dina = {96'd0, 16'd33350, 16'd36472, 16'd43947, 16'd27480, 16'd64400, 16'd6289, 16'd10575, 16'd16156, 16'd48577, 16'd50680}; // indx = 999
    #10;
    addra = 32'd32000;
    dina = {96'd0, 16'd2698, 16'd56115, 16'd20164, 16'd880, 16'd40757, 16'd15467, 16'd18017, 16'd63382, 16'd46378, 16'd45776}; // indx = 1000
    #10;
    addra = 32'd32032;
    dina = {96'd0, 16'd39193, 16'd27076, 16'd35756, 16'd31378, 16'd21132, 16'd14342, 16'd28282, 16'd22097, 16'd5487, 16'd5210}; // indx = 1001
    #10;
    addra = 32'd32064;
    dina = {96'd0, 16'd57015, 16'd14163, 16'd52751, 16'd20898, 16'd16003, 16'd14691, 16'd35935, 16'd3635, 16'd44797, 16'd24240}; // indx = 1002
    #10;
    addra = 32'd32096;
    dina = {96'd0, 16'd62056, 16'd38789, 16'd47880, 16'd7157, 16'd2755, 16'd45682, 16'd45763, 16'd26369, 16'd4346, 16'd15589}; // indx = 1003
    #10;
    addra = 32'd32128;
    dina = {96'd0, 16'd27928, 16'd56548, 16'd22292, 16'd61165, 16'd34932, 16'd845, 16'd35066, 16'd18497, 16'd322, 16'd27552}; // indx = 1004
    #10;
    addra = 32'd32160;
    dina = {96'd0, 16'd41058, 16'd1023, 16'd6305, 16'd60566, 16'd17228, 16'd36281, 16'd26, 16'd39714, 16'd44694, 16'd60892}; // indx = 1005
    #10;
    addra = 32'd32192;
    dina = {96'd0, 16'd51515, 16'd39629, 16'd18518, 16'd24517, 16'd63984, 16'd54362, 16'd42903, 16'd58897, 16'd10668, 16'd8411}; // indx = 1006
    #10;
    addra = 32'd32224;
    dina = {96'd0, 16'd63297, 16'd13894, 16'd52545, 16'd5298, 16'd29473, 16'd42315, 16'd36875, 16'd46455, 16'd59298, 16'd1626}; // indx = 1007
    #10;
    addra = 32'd32256;
    dina = {96'd0, 16'd12948, 16'd39879, 16'd20190, 16'd48897, 16'd49319, 16'd45940, 16'd27919, 16'd24344, 16'd45154, 16'd17975}; // indx = 1008
    #10;
    addra = 32'd32288;
    dina = {96'd0, 16'd27363, 16'd16468, 16'd56830, 16'd50587, 16'd53771, 16'd49693, 16'd48182, 16'd3948, 16'd39372, 16'd38849}; // indx = 1009
    #10;
    addra = 32'd32320;
    dina = {96'd0, 16'd15408, 16'd35201, 16'd22337, 16'd10176, 16'd35518, 16'd58800, 16'd5595, 16'd23554, 16'd30816, 16'd61322}; // indx = 1010
    #10;
    addra = 32'd32352;
    dina = {96'd0, 16'd44882, 16'd33250, 16'd461, 16'd32298, 16'd55572, 16'd23127, 16'd16519, 16'd51047, 16'd56135, 16'd54167}; // indx = 1011
    #10;
    addra = 32'd32384;
    dina = {96'd0, 16'd49907, 16'd55866, 16'd25155, 16'd62267, 16'd29099, 16'd16777, 16'd17826, 16'd9161, 16'd25848, 16'd57855}; // indx = 1012
    #10;
    addra = 32'd32416;
    dina = {96'd0, 16'd42703, 16'd4448, 16'd34723, 16'd29201, 16'd31901, 16'd8224, 16'd48941, 16'd35584, 16'd50189, 16'd15215}; // indx = 1013
    #10;
    addra = 32'd32448;
    dina = {96'd0, 16'd17509, 16'd15734, 16'd17305, 16'd36985, 16'd58306, 16'd43243, 16'd43908, 16'd26181, 16'd17887, 16'd40313}; // indx = 1014
    #10;
    addra = 32'd32480;
    dina = {96'd0, 16'd62782, 16'd9505, 16'd48871, 16'd13076, 16'd25490, 16'd20699, 16'd34550, 16'd2448, 16'd26270, 16'd6717}; // indx = 1015
    #10;
    addra = 32'd32512;
    dina = {96'd0, 16'd56864, 16'd31097, 16'd17699, 16'd46360, 16'd35190, 16'd29374, 16'd64292, 16'd20394, 16'd52282, 16'd47459}; // indx = 1016
    #10;
    addra = 32'd32544;
    dina = {96'd0, 16'd61393, 16'd17528, 16'd26946, 16'd62217, 16'd55792, 16'd41940, 16'd18309, 16'd63398, 16'd7647, 16'd55525}; // indx = 1017
    #10;
    addra = 32'd32576;
    dina = {96'd0, 16'd11837, 16'd51654, 16'd56698, 16'd52065, 16'd14736, 16'd20906, 16'd4295, 16'd38895, 16'd23256, 16'd35043}; // indx = 1018
    #10;
    addra = 32'd32608;
    dina = {96'd0, 16'd55527, 16'd1354, 16'd30483, 16'd15804, 16'd34416, 16'd45072, 16'd31493, 16'd27095, 16'd40280, 16'd10374}; // indx = 1019
    #10;
    addra = 32'd32640;
    dina = {96'd0, 16'd4614, 16'd43078, 16'd39232, 16'd1462, 16'd50358, 16'd39911, 16'd28697, 16'd41664, 16'd62171, 16'd2638}; // indx = 1020
    #10;
    addra = 32'd32672;
    dina = {96'd0, 16'd32846, 16'd57153, 16'd44326, 16'd60431, 16'd50808, 16'd16756, 16'd50300, 16'd7094, 16'd37139, 16'd9750}; // indx = 1021
    #10;
    addra = 32'd32704;
    dina = {96'd0, 16'd763, 16'd46693, 16'd38791, 16'd4808, 16'd18300, 16'd6227, 16'd23377, 16'd12579, 16'd34292, 16'd43274}; // indx = 1022
    #10;
    addra = 32'd32736;
    dina = {96'd0, 16'd52382, 16'd4396, 16'd15971, 16'd18967, 16'd27354, 16'd47775, 16'd36874, 16'd32744, 16'd30904, 16'd4611}; // indx = 1023
    #10;
    addra = 32'd32768;
    dina = {96'd0, 16'd4973, 16'd49860, 16'd13243, 16'd41796, 16'd23822, 16'd26302, 16'd9210, 16'd35795, 16'd18814, 16'd41223}; // indx = 1024
    #10;
    addra = 32'd32800;
    dina = {96'd0, 16'd39531, 16'd21370, 16'd12969, 16'd46369, 16'd10666, 16'd64111, 16'd47445, 16'd62245, 16'd32444, 16'd2991}; // indx = 1025
    #10;
    addra = 32'd32832;
    dina = {96'd0, 16'd37549, 16'd56974, 16'd51138, 16'd20240, 16'd54154, 16'd5693, 16'd3305, 16'd10211, 16'd58091, 16'd14354}; // indx = 1026
    #10;
    addra = 32'd32864;
    dina = {96'd0, 16'd39064, 16'd13326, 16'd11577, 16'd24439, 16'd41885, 16'd19714, 16'd45457, 16'd51473, 16'd56945, 16'd26090}; // indx = 1027
    #10;
    addra = 32'd32896;
    dina = {96'd0, 16'd54989, 16'd42626, 16'd1741, 16'd37912, 16'd20485, 16'd191, 16'd14069, 16'd13436, 16'd9315, 16'd61113}; // indx = 1028
    #10;
    addra = 32'd32928;
    dina = {96'd0, 16'd42386, 16'd19389, 16'd29550, 16'd61626, 16'd18929, 16'd11714, 16'd10583, 16'd4883, 16'd60313, 16'd8322}; // indx = 1029
    #10;
    addra = 32'd32960;
    dina = {96'd0, 16'd63835, 16'd15191, 16'd8891, 16'd9061, 16'd34847, 16'd28172, 16'd57301, 16'd35899, 16'd59392, 16'd47602}; // indx = 1030
    #10;
    addra = 32'd32992;
    dina = {96'd0, 16'd41172, 16'd11928, 16'd30293, 16'd50567, 16'd41754, 16'd62123, 16'd6546, 16'd10286, 16'd64480, 16'd24238}; // indx = 1031
    #10;
    addra = 32'd33024;
    dina = {96'd0, 16'd15269, 16'd37784, 16'd3915, 16'd23297, 16'd62665, 16'd47618, 16'd48874, 16'd782, 16'd34698, 16'd65032}; // indx = 1032
    #10;
    addra = 32'd33056;
    dina = {96'd0, 16'd39298, 16'd25556, 16'd7592, 16'd38022, 16'd52806, 16'd5425, 16'd2900, 16'd11324, 16'd52818, 16'd32879}; // indx = 1033
    #10;
    addra = 32'd33088;
    dina = {96'd0, 16'd43989, 16'd49122, 16'd44992, 16'd37209, 16'd40328, 16'd1348, 16'd23836, 16'd13127, 16'd14869, 16'd57288}; // indx = 1034
    #10;
    addra = 32'd33120;
    dina = {96'd0, 16'd21781, 16'd19654, 16'd29149, 16'd5525, 16'd27375, 16'd12947, 16'd33355, 16'd26007, 16'd23512, 16'd64439}; // indx = 1035
    #10;
    addra = 32'd33152;
    dina = {96'd0, 16'd15812, 16'd30011, 16'd47273, 16'd29038, 16'd17044, 16'd64033, 16'd32058, 16'd65104, 16'd30811, 16'd58151}; // indx = 1036
    #10;
    addra = 32'd33184;
    dina = {96'd0, 16'd36229, 16'd6065, 16'd31249, 16'd56488, 16'd38131, 16'd46228, 16'd8350, 16'd38620, 16'd20721, 16'd6704}; // indx = 1037
    #10;
    addra = 32'd33216;
    dina = {96'd0, 16'd48048, 16'd15451, 16'd25166, 16'd10924, 16'd15232, 16'd29910, 16'd51146, 16'd13970, 16'd56323, 16'd12424}; // indx = 1038
    #10;
    addra = 32'd33248;
    dina = {96'd0, 16'd11157, 16'd13588, 16'd42044, 16'd64314, 16'd4243, 16'd12448, 16'd51483, 16'd60768, 16'd47435, 16'd63804}; // indx = 1039
    #10;
    addra = 32'd33280;
    dina = {96'd0, 16'd54984, 16'd40682, 16'd7678, 16'd54381, 16'd32460, 16'd37560, 16'd20366, 16'd62722, 16'd39609, 16'd59894}; // indx = 1040
    #10;
    addra = 32'd33312;
    dina = {96'd0, 16'd32264, 16'd58328, 16'd50298, 16'd27310, 16'd52493, 16'd49201, 16'd47818, 16'd11012, 16'd3931, 16'd4736}; // indx = 1041
    #10;
    addra = 32'd33344;
    dina = {96'd0, 16'd46533, 16'd13186, 16'd34179, 16'd6115, 16'd60779, 16'd33490, 16'd16296, 16'd12704, 16'd56586, 16'd23145}; // indx = 1042
    #10;
    addra = 32'd33376;
    dina = {96'd0, 16'd32637, 16'd35478, 16'd28943, 16'd5655, 16'd58428, 16'd39395, 16'd24048, 16'd12119, 16'd21029, 16'd39115}; // indx = 1043
    #10;
    addra = 32'd33408;
    dina = {96'd0, 16'd11075, 16'd33472, 16'd52521, 16'd20535, 16'd20264, 16'd20583, 16'd44026, 16'd37078, 16'd51942, 16'd49389}; // indx = 1044
    #10;
    addra = 32'd33440;
    dina = {96'd0, 16'd2768, 16'd2643, 16'd26274, 16'd3064, 16'd679, 16'd42507, 16'd41486, 16'd60909, 16'd4995, 16'd40334}; // indx = 1045
    #10;
    addra = 32'd33472;
    dina = {96'd0, 16'd39523, 16'd2836, 16'd56592, 16'd2947, 16'd41586, 16'd29647, 16'd35150, 16'd4696, 16'd55746, 16'd49820}; // indx = 1046
    #10;
    addra = 32'd33504;
    dina = {96'd0, 16'd45509, 16'd24691, 16'd65263, 16'd51156, 16'd61389, 16'd16861, 16'd20712, 16'd13665, 16'd27315, 16'd44956}; // indx = 1047
    #10;
    addra = 32'd33536;
    dina = {96'd0, 16'd64646, 16'd61044, 16'd41351, 16'd60538, 16'd43058, 16'd61734, 16'd47740, 16'd42121, 16'd46975, 16'd42619}; // indx = 1048
    #10;
    addra = 32'd33568;
    dina = {96'd0, 16'd6926, 16'd9399, 16'd44942, 16'd25969, 16'd28950, 16'd57227, 16'd28758, 16'd56611, 16'd47859, 16'd28975}; // indx = 1049
    #10;
    addra = 32'd33600;
    dina = {96'd0, 16'd28186, 16'd46575, 16'd21770, 16'd15090, 16'd41861, 16'd36852, 16'd21363, 16'd33442, 16'd1790, 16'd27733}; // indx = 1050
    #10;
    addra = 32'd33632;
    dina = {96'd0, 16'd36637, 16'd23224, 16'd64945, 16'd26367, 16'd52518, 16'd10904, 16'd32765, 16'd547, 16'd11631, 16'd33324}; // indx = 1051
    #10;
    addra = 32'd33664;
    dina = {96'd0, 16'd5039, 16'd25473, 16'd44272, 16'd6919, 16'd49271, 16'd49603, 16'd54469, 16'd3048, 16'd56107, 16'd50692}; // indx = 1052
    #10;
    addra = 32'd33696;
    dina = {96'd0, 16'd17763, 16'd18569, 16'd24971, 16'd31894, 16'd3556, 16'd12118, 16'd46072, 16'd47380, 16'd6807, 16'd44282}; // indx = 1053
    #10;
    addra = 32'd33728;
    dina = {96'd0, 16'd12857, 16'd64293, 16'd14326, 16'd61755, 16'd3342, 16'd13747, 16'd21195, 16'd15926, 16'd62247, 16'd49618}; // indx = 1054
    #10;
    addra = 32'd33760;
    dina = {96'd0, 16'd17612, 16'd37919, 16'd27733, 16'd14827, 16'd22004, 16'd57820, 16'd55034, 16'd53593, 16'd57832, 16'd23185}; // indx = 1055
    #10;
    addra = 32'd33792;
    dina = {96'd0, 16'd37237, 16'd5641, 16'd1491, 16'd7816, 16'd59961, 16'd63339, 16'd42474, 16'd35594, 16'd7613, 16'd3983}; // indx = 1056
    #10;
    addra = 32'd33824;
    dina = {96'd0, 16'd34338, 16'd10808, 16'd19386, 16'd61422, 16'd57395, 16'd2538, 16'd43132, 16'd29899, 16'd61819, 16'd35394}; // indx = 1057
    #10;
    addra = 32'd33856;
    dina = {96'd0, 16'd27211, 16'd55984, 16'd32181, 16'd19533, 16'd2920, 16'd1371, 16'd41408, 16'd11342, 16'd37361, 16'd866}; // indx = 1058
    #10;
    addra = 32'd33888;
    dina = {96'd0, 16'd46247, 16'd19649, 16'd56222, 16'd49806, 16'd57061, 16'd18611, 16'd56128, 16'd61132, 16'd20326, 16'd56452}; // indx = 1059
    #10;
    addra = 32'd33920;
    dina = {96'd0, 16'd20457, 16'd17988, 16'd8067, 16'd26862, 16'd20831, 16'd57884, 16'd12042, 16'd43785, 16'd61299, 16'd44262}; // indx = 1060
    #10;
    addra = 32'd33952;
    dina = {96'd0, 16'd37128, 16'd8829, 16'd60698, 16'd23935, 16'd47024, 16'd7728, 16'd4073, 16'd52238, 16'd27217, 16'd41510}; // indx = 1061
    #10;
    addra = 32'd33984;
    dina = {96'd0, 16'd46089, 16'd42316, 16'd12451, 16'd23396, 16'd24890, 16'd25478, 16'd57324, 16'd51576, 16'd24413, 16'd9306}; // indx = 1062
    #10;
    addra = 32'd34016;
    dina = {96'd0, 16'd6726, 16'd46158, 16'd1414, 16'd8055, 16'd6621, 16'd30679, 16'd46888, 16'd32137, 16'd446, 16'd62977}; // indx = 1063
    #10;
    addra = 32'd34048;
    dina = {96'd0, 16'd51594, 16'd34026, 16'd55359, 16'd33178, 16'd45854, 16'd52493, 16'd8473, 16'd6118, 16'd649, 16'd38207}; // indx = 1064
    #10;
    addra = 32'd34080;
    dina = {96'd0, 16'd3526, 16'd14017, 16'd61952, 16'd15984, 16'd58818, 16'd50411, 16'd15847, 16'd57591, 16'd13190, 16'd21074}; // indx = 1065
    #10;
    addra = 32'd34112;
    dina = {96'd0, 16'd48434, 16'd51509, 16'd21028, 16'd57498, 16'd10315, 16'd11592, 16'd45361, 16'd64985, 16'd23157, 16'd63677}; // indx = 1066
    #10;
    addra = 32'd34144;
    dina = {96'd0, 16'd64133, 16'd60991, 16'd33204, 16'd42576, 16'd6348, 16'd1383, 16'd42187, 16'd32021, 16'd32622, 16'd51704}; // indx = 1067
    #10;
    addra = 32'd34176;
    dina = {96'd0, 16'd2451, 16'd18912, 16'd27754, 16'd22448, 16'd42003, 16'd6958, 16'd7863, 16'd63897, 16'd16038, 16'd9967}; // indx = 1068
    #10;
    addra = 32'd34208;
    dina = {96'd0, 16'd49643, 16'd33999, 16'd52761, 16'd4034, 16'd6992, 16'd46049, 16'd2563, 16'd814, 16'd26459, 16'd28381}; // indx = 1069
    #10;
    addra = 32'd34240;
    dina = {96'd0, 16'd25377, 16'd15091, 16'd35172, 16'd10084, 16'd47095, 16'd31673, 16'd64078, 16'd725, 16'd14408, 16'd33064}; // indx = 1070
    #10;
    addra = 32'd34272;
    dina = {96'd0, 16'd27298, 16'd64334, 16'd38558, 16'd39997, 16'd26426, 16'd31543, 16'd44720, 16'd56692, 16'd42292, 16'd59141}; // indx = 1071
    #10;
    addra = 32'd34304;
    dina = {96'd0, 16'd36910, 16'd58870, 16'd38217, 16'd26175, 16'd44136, 16'd58811, 16'd50930, 16'd64211, 16'd63200, 16'd12751}; // indx = 1072
    #10;
    addra = 32'd34336;
    dina = {96'd0, 16'd16981, 16'd54461, 16'd35151, 16'd46894, 16'd53563, 16'd33746, 16'd26801, 16'd34443, 16'd52563, 16'd54656}; // indx = 1073
    #10;
    addra = 32'd34368;
    dina = {96'd0, 16'd33801, 16'd8012, 16'd22255, 16'd47473, 16'd58630, 16'd9943, 16'd16257, 16'd31994, 16'd971, 16'd27891}; // indx = 1074
    #10;
    addra = 32'd34400;
    dina = {96'd0, 16'd64353, 16'd12094, 16'd43654, 16'd4231, 16'd33603, 16'd6193, 16'd49449, 16'd50339, 16'd43386, 16'd53856}; // indx = 1075
    #10;
    addra = 32'd34432;
    dina = {96'd0, 16'd58220, 16'd39389, 16'd24106, 16'd21703, 16'd64450, 16'd36888, 16'd17318, 16'd50478, 16'd31239, 16'd41864}; // indx = 1076
    #10;
    addra = 32'd34464;
    dina = {96'd0, 16'd48630, 16'd48430, 16'd48830, 16'd40497, 16'd38519, 16'd27516, 16'd40134, 16'd31691, 16'd20456, 16'd63353}; // indx = 1077
    #10;
    addra = 32'd34496;
    dina = {96'd0, 16'd46172, 16'd8945, 16'd28474, 16'd33602, 16'd47962, 16'd19361, 16'd21909, 16'd742, 16'd46459, 16'd24855}; // indx = 1078
    #10;
    addra = 32'd34528;
    dina = {96'd0, 16'd41516, 16'd54075, 16'd10099, 16'd31555, 16'd15812, 16'd16711, 16'd51177, 16'd57042, 16'd19113, 16'd32660}; // indx = 1079
    #10;
    addra = 32'd34560;
    dina = {96'd0, 16'd23918, 16'd48175, 16'd58696, 16'd50074, 16'd53052, 16'd61099, 16'd12509, 16'd9177, 16'd31623, 16'd18355}; // indx = 1080
    #10;
    addra = 32'd34592;
    dina = {96'd0, 16'd28306, 16'd55874, 16'd11422, 16'd44705, 16'd25528, 16'd21996, 16'd34149, 16'd30453, 16'd11481, 16'd7909}; // indx = 1081
    #10;
    addra = 32'd34624;
    dina = {96'd0, 16'd55807, 16'd2441, 16'd48483, 16'd30859, 16'd9180, 16'd40625, 16'd3082, 16'd19024, 16'd4791, 16'd38048}; // indx = 1082
    #10;
    addra = 32'd34656;
    dina = {96'd0, 16'd43398, 16'd1238, 16'd38920, 16'd25853, 16'd53744, 16'd5604, 16'd60167, 16'd56500, 16'd56216, 16'd222}; // indx = 1083
    #10;
    addra = 32'd34688;
    dina = {96'd0, 16'd1851, 16'd48202, 16'd31922, 16'd28314, 16'd56446, 16'd38715, 16'd31313, 16'd9282, 16'd7132, 16'd12076}; // indx = 1084
    #10;
    addra = 32'd34720;
    dina = {96'd0, 16'd47090, 16'd59854, 16'd11181, 16'd54149, 16'd60474, 16'd54823, 16'd28301, 16'd62567, 16'd24688, 16'd61488}; // indx = 1085
    #10;
    addra = 32'd34752;
    dina = {96'd0, 16'd21700, 16'd107, 16'd40318, 16'd15083, 16'd60444, 16'd3775, 16'd9967, 16'd23348, 16'd56155, 16'd19782}; // indx = 1086
    #10;
    addra = 32'd34784;
    dina = {96'd0, 16'd17036, 16'd64834, 16'd45490, 16'd12567, 16'd7696, 16'd926, 16'd48626, 16'd2528, 16'd40195, 16'd4329}; // indx = 1087
    #10;
    addra = 32'd34816;
    dina = {96'd0, 16'd20587, 16'd18188, 16'd59367, 16'd10720, 16'd24568, 16'd27974, 16'd10260, 16'd62073, 16'd24226, 16'd59777}; // indx = 1088
    #10;
    addra = 32'd34848;
    dina = {96'd0, 16'd28995, 16'd39693, 16'd44859, 16'd40203, 16'd50582, 16'd61758, 16'd20295, 16'd12729, 16'd33410, 16'd13019}; // indx = 1089
    #10;
    addra = 32'd34880;
    dina = {96'd0, 16'd50144, 16'd39708, 16'd10269, 16'd44236, 16'd39838, 16'd28094, 16'd6070, 16'd38580, 16'd39892, 16'd24388}; // indx = 1090
    #10;
    addra = 32'd34912;
    dina = {96'd0, 16'd33385, 16'd64966, 16'd18818, 16'd13885, 16'd65221, 16'd9158, 16'd21645, 16'd25361, 16'd24181, 16'd55239}; // indx = 1091
    #10;
    addra = 32'd34944;
    dina = {96'd0, 16'd13958, 16'd39951, 16'd12593, 16'd20240, 16'd25961, 16'd1347, 16'd33828, 16'd57609, 16'd39305, 16'd27929}; // indx = 1092
    #10;
    addra = 32'd34976;
    dina = {96'd0, 16'd30198, 16'd25722, 16'd33021, 16'd42972, 16'd25437, 16'd2344, 16'd65179, 16'd59766, 16'd58722, 16'd48660}; // indx = 1093
    #10;
    addra = 32'd35008;
    dina = {96'd0, 16'd18329, 16'd27777, 16'd21779, 16'd12518, 16'd20284, 16'd38887, 16'd21408, 16'd57438, 16'd60870, 16'd43257}; // indx = 1094
    #10;
    addra = 32'd35040;
    dina = {96'd0, 16'd16371, 16'd30274, 16'd31435, 16'd38715, 16'd33364, 16'd8760, 16'd41596, 16'd55663, 16'd29609, 16'd13657}; // indx = 1095
    #10;
    addra = 32'd35072;
    dina = {96'd0, 16'd61790, 16'd52739, 16'd2881, 16'd29871, 16'd39542, 16'd48678, 16'd47537, 16'd31347, 16'd5203, 16'd48035}; // indx = 1096
    #10;
    addra = 32'd35104;
    dina = {96'd0, 16'd17436, 16'd17162, 16'd53260, 16'd50268, 16'd42452, 16'd31269, 16'd62417, 16'd32578, 16'd36800, 16'd11999}; // indx = 1097
    #10;
    addra = 32'd35136;
    dina = {96'd0, 16'd14412, 16'd51211, 16'd20936, 16'd4861, 16'd27973, 16'd46696, 16'd58589, 16'd21016, 16'd45640, 16'd53643}; // indx = 1098
    #10;
    addra = 32'd35168;
    dina = {96'd0, 16'd24681, 16'd20682, 16'd14585, 16'd30589, 16'd205, 16'd39801, 16'd1227, 16'd22215, 16'd58027, 16'd52479}; // indx = 1099
    #10;
    addra = 32'd35200;
    dina = {96'd0, 16'd18845, 16'd17288, 16'd39134, 16'd45025, 16'd62800, 16'd56655, 16'd37749, 16'd30378, 16'd38942, 16'd44310}; // indx = 1100
    #10;
    addra = 32'd35232;
    dina = {96'd0, 16'd35939, 16'd56643, 16'd44350, 16'd48324, 16'd51666, 16'd19521, 16'd41930, 16'd30724, 16'd39445, 16'd29453}; // indx = 1101
    #10;
    addra = 32'd35264;
    dina = {96'd0, 16'd42911, 16'd43818, 16'd13593, 16'd59548, 16'd12506, 16'd31890, 16'd12615, 16'd13232, 16'd29325, 16'd40343}; // indx = 1102
    #10;
    addra = 32'd35296;
    dina = {96'd0, 16'd12178, 16'd62373, 16'd17964, 16'd8863, 16'd14454, 16'd23150, 16'd7214, 16'd891, 16'd48300, 16'd8593}; // indx = 1103
    #10;
    addra = 32'd35328;
    dina = {96'd0, 16'd243, 16'd63232, 16'd61886, 16'd26697, 16'd18800, 16'd533, 16'd11775, 16'd35112, 16'd36387, 16'd24117}; // indx = 1104
    #10;
    addra = 32'd35360;
    dina = {96'd0, 16'd27033, 16'd23919, 16'd56253, 16'd25898, 16'd8463, 16'd12150, 16'd63594, 16'd30841, 16'd2091, 16'd64335}; // indx = 1105
    #10;
    addra = 32'd35392;
    dina = {96'd0, 16'd54685, 16'd41449, 16'd13433, 16'd13462, 16'd14895, 16'd65450, 16'd30942, 16'd19715, 16'd62460, 16'd54217}; // indx = 1106
    #10;
    addra = 32'd35424;
    dina = {96'd0, 16'd12347, 16'd35660, 16'd49000, 16'd15656, 16'd2416, 16'd46196, 16'd43264, 16'd21286, 16'd9331, 16'd41635}; // indx = 1107
    #10;
    addra = 32'd35456;
    dina = {96'd0, 16'd59192, 16'd64627, 16'd16643, 16'd54464, 16'd41131, 16'd8427, 16'd21942, 16'd19394, 16'd31573, 16'd40658}; // indx = 1108
    #10;
    addra = 32'd35488;
    dina = {96'd0, 16'd7127, 16'd43389, 16'd34039, 16'd60809, 16'd38813, 16'd63624, 16'd57605, 16'd15695, 16'd26705, 16'd29762}; // indx = 1109
    #10;
    addra = 32'd35520;
    dina = {96'd0, 16'd29507, 16'd3246, 16'd1689, 16'd39336, 16'd53623, 16'd54899, 16'd25170, 16'd35109, 16'd524, 16'd41324}; // indx = 1110
    #10;
    addra = 32'd35552;
    dina = {96'd0, 16'd5573, 16'd11887, 16'd63050, 16'd46984, 16'd28870, 16'd36831, 16'd57436, 16'd50059, 16'd4224, 16'd54006}; // indx = 1111
    #10;
    addra = 32'd35584;
    dina = {96'd0, 16'd8654, 16'd54218, 16'd22912, 16'd62422, 16'd10437, 16'd59302, 16'd45091, 16'd17284, 16'd52542, 16'd11244}; // indx = 1112
    #10;
    addra = 32'd35616;
    dina = {96'd0, 16'd3694, 16'd37877, 16'd4214, 16'd18328, 16'd22512, 16'd23171, 16'd34575, 16'd58097, 16'd32760, 16'd17953}; // indx = 1113
    #10;
    addra = 32'd35648;
    dina = {96'd0, 16'd2511, 16'd661, 16'd38401, 16'd7554, 16'd51281, 16'd60671, 16'd35272, 16'd40443, 16'd61283, 16'd11812}; // indx = 1114
    #10;
    addra = 32'd35680;
    dina = {96'd0, 16'd30992, 16'd49715, 16'd30220, 16'd2563, 16'd35314, 16'd53820, 16'd13418, 16'd56896, 16'd32373, 16'd1526}; // indx = 1115
    #10;
    addra = 32'd35712;
    dina = {96'd0, 16'd2494, 16'd15824, 16'd18066, 16'd50798, 16'd19341, 16'd64946, 16'd16632, 16'd48409, 16'd42728, 16'd21314}; // indx = 1116
    #10;
    addra = 32'd35744;
    dina = {96'd0, 16'd49232, 16'd18398, 16'd16972, 16'd64872, 16'd15572, 16'd47123, 16'd31217, 16'd24468, 16'd36018, 16'd28669}; // indx = 1117
    #10;
    addra = 32'd35776;
    dina = {96'd0, 16'd392, 16'd47612, 16'd64217, 16'd9354, 16'd57201, 16'd48081, 16'd19785, 16'd40206, 16'd5027, 16'd40440}; // indx = 1118
    #10;
    addra = 32'd35808;
    dina = {96'd0, 16'd62634, 16'd25639, 16'd2501, 16'd3192, 16'd24076, 16'd24328, 16'd34070, 16'd42454, 16'd6056, 16'd24571}; // indx = 1119
    #10;
    addra = 32'd35840;
    dina = {96'd0, 16'd50944, 16'd53740, 16'd20576, 16'd62733, 16'd23999, 16'd30149, 16'd1917, 16'd3438, 16'd64784, 16'd41361}; // indx = 1120
    #10;
    addra = 32'd35872;
    dina = {96'd0, 16'd47908, 16'd59984, 16'd61938, 16'd49762, 16'd20437, 16'd6925, 16'd11565, 16'd51548, 16'd13792, 16'd63150}; // indx = 1121
    #10;
    addra = 32'd35904;
    dina = {96'd0, 16'd36918, 16'd57743, 16'd18786, 16'd19297, 16'd54591, 16'd37489, 16'd2887, 16'd50024, 16'd2324, 16'd5520}; // indx = 1122
    #10;
    addra = 32'd35936;
    dina = {96'd0, 16'd47723, 16'd23670, 16'd54597, 16'd20733, 16'd28677, 16'd46888, 16'd41544, 16'd2670, 16'd12785, 16'd47370}; // indx = 1123
    #10;
    addra = 32'd35968;
    dina = {96'd0, 16'd54791, 16'd18161, 16'd16904, 16'd19907, 16'd1905, 16'd57517, 16'd28284, 16'd9023, 16'd56586, 16'd16789}; // indx = 1124
    #10;
    addra = 32'd36000;
    dina = {96'd0, 16'd7702, 16'd61247, 16'd64854, 16'd15967, 16'd44077, 16'd24312, 16'd58945, 16'd46545, 16'd4174, 16'd8919}; // indx = 1125
    #10;
    addra = 32'd36032;
    dina = {96'd0, 16'd32022, 16'd9522, 16'd20942, 16'd49712, 16'd1342, 16'd2769, 16'd52449, 16'd2010, 16'd31581, 16'd511}; // indx = 1126
    #10;
    addra = 32'd36064;
    dina = {96'd0, 16'd34969, 16'd51399, 16'd38214, 16'd37770, 16'd43035, 16'd13398, 16'd47353, 16'd49141, 16'd43039, 16'd16220}; // indx = 1127
    #10;
    addra = 32'd36096;
    dina = {96'd0, 16'd8096, 16'd63799, 16'd7633, 16'd3473, 16'd41030, 16'd18810, 16'd56516, 16'd31033, 16'd27, 16'd53273}; // indx = 1128
    #10;
    addra = 32'd36128;
    dina = {96'd0, 16'd41238, 16'd4682, 16'd3083, 16'd42248, 16'd21662, 16'd31570, 16'd50823, 16'd24710, 16'd22437, 16'd60030}; // indx = 1129
    #10;
    addra = 32'd36160;
    dina = {96'd0, 16'd57382, 16'd52516, 16'd44322, 16'd43381, 16'd44788, 16'd60889, 16'd29828, 16'd24272, 16'd62757, 16'd37068}; // indx = 1130
    #10;
    addra = 32'd36192;
    dina = {96'd0, 16'd48487, 16'd18176, 16'd27334, 16'd11265, 16'd54924, 16'd2363, 16'd23264, 16'd58235, 16'd8466, 16'd57}; // indx = 1131
    #10;
    addra = 32'd36224;
    dina = {96'd0, 16'd25065, 16'd17031, 16'd60266, 16'd1476, 16'd5037, 16'd40224, 16'd43676, 16'd32162, 16'd8467, 16'd34876}; // indx = 1132
    #10;
    addra = 32'd36256;
    dina = {96'd0, 16'd16236, 16'd9243, 16'd6270, 16'd33204, 16'd6450, 16'd5949, 16'd19653, 16'd5306, 16'd17472, 16'd27355}; // indx = 1133
    #10;
    addra = 32'd36288;
    dina = {96'd0, 16'd17532, 16'd13711, 16'd53103, 16'd6405, 16'd14655, 16'd34734, 16'd11664, 16'd34044, 16'd28369, 16'd7056}; // indx = 1134
    #10;
    addra = 32'd36320;
    dina = {96'd0, 16'd17516, 16'd63188, 16'd11294, 16'd15697, 16'd3652, 16'd50050, 16'd62859, 16'd5252, 16'd57916, 16'd58801}; // indx = 1135
    #10;
    addra = 32'd36352;
    dina = {96'd0, 16'd64352, 16'd23654, 16'd973, 16'd11823, 16'd54353, 16'd2843, 16'd59964, 16'd55178, 16'd27356, 16'd3537}; // indx = 1136
    #10;
    addra = 32'd36384;
    dina = {96'd0, 16'd8114, 16'd771, 16'd40057, 16'd17659, 16'd64060, 16'd22686, 16'd59006, 16'd28845, 16'd15850, 16'd6386}; // indx = 1137
    #10;
    addra = 32'd36416;
    dina = {96'd0, 16'd32317, 16'd10029, 16'd3174, 16'd34538, 16'd2485, 16'd57984, 16'd47573, 16'd48667, 16'd1265, 16'd34946}; // indx = 1138
    #10;
    addra = 32'd36448;
    dina = {96'd0, 16'd15580, 16'd16538, 16'd33666, 16'd64608, 16'd13225, 16'd44380, 16'd17006, 16'd39723, 16'd28272, 16'd13800}; // indx = 1139
    #10;
    addra = 32'd36480;
    dina = {96'd0, 16'd54414, 16'd20596, 16'd33728, 16'd62765, 16'd34068, 16'd48941, 16'd42234, 16'd56491, 16'd23517, 16'd29483}; // indx = 1140
    #10;
    addra = 32'd36512;
    dina = {96'd0, 16'd59904, 16'd29417, 16'd10650, 16'd7122, 16'd14627, 16'd43064, 16'd57246, 16'd9874, 16'd63305, 16'd11941}; // indx = 1141
    #10;
    addra = 32'd36544;
    dina = {96'd0, 16'd18901, 16'd64161, 16'd2876, 16'd33745, 16'd9975, 16'd21729, 16'd25803, 16'd10419, 16'd47645, 16'd30272}; // indx = 1142
    #10;
    addra = 32'd36576;
    dina = {96'd0, 16'd30881, 16'd60870, 16'd25091, 16'd58592, 16'd21587, 16'd50881, 16'd14081, 16'd12594, 16'd63943, 16'd54196}; // indx = 1143
    #10;
    addra = 32'd36608;
    dina = {96'd0, 16'd17136, 16'd20251, 16'd41933, 16'd42842, 16'd12050, 16'd12811, 16'd3933, 16'd61542, 16'd38559, 16'd54049}; // indx = 1144
    #10;
    addra = 32'd36640;
    dina = {96'd0, 16'd14004, 16'd45955, 16'd27482, 16'd47429, 16'd20434, 16'd9126, 16'd7438, 16'd58451, 16'd58312, 16'd4345}; // indx = 1145
    #10;
    addra = 32'd36672;
    dina = {96'd0, 16'd27906, 16'd16870, 16'd39391, 16'd12845, 16'd24357, 16'd32455, 16'd22844, 16'd18612, 16'd58833, 16'd51201}; // indx = 1146
    #10;
    addra = 32'd36704;
    dina = {96'd0, 16'd40317, 16'd14044, 16'd26060, 16'd12205, 16'd20229, 16'd23762, 16'd51573, 16'd2608, 16'd23409, 16'd8859}; // indx = 1147
    #10;
    addra = 32'd36736;
    dina = {96'd0, 16'd2049, 16'd38120, 16'd20031, 16'd58917, 16'd42121, 16'd25316, 16'd27445, 16'd5940, 16'd24136, 16'd65413}; // indx = 1148
    #10;
    addra = 32'd36768;
    dina = {96'd0, 16'd17396, 16'd11259, 16'd28822, 16'd9388, 16'd19385, 16'd35528, 16'd18391, 16'd13688, 16'd38740, 16'd52440}; // indx = 1149
    #10;
    addra = 32'd36800;
    dina = {96'd0, 16'd22568, 16'd33118, 16'd20188, 16'd16450, 16'd41947, 16'd33455, 16'd63962, 16'd2688, 16'd52736, 16'd61453}; // indx = 1150
    #10;
    addra = 32'd36832;
    dina = {96'd0, 16'd6169, 16'd15343, 16'd48962, 16'd52205, 16'd20305, 16'd65513, 16'd36125, 16'd65065, 16'd12631, 16'd4910}; // indx = 1151
    #10;
    addra = 32'd36864;
    dina = {96'd0, 16'd9033, 16'd25235, 16'd52513, 16'd46449, 16'd52287, 16'd46296, 16'd53224, 16'd32629, 16'd33136, 16'd39563}; // indx = 1152
    #10;
    addra = 32'd36896;
    dina = {96'd0, 16'd1703, 16'd62593, 16'd52823, 16'd11343, 16'd5688, 16'd17845, 16'd58054, 16'd57518, 16'd49869, 16'd47593}; // indx = 1153
    #10;
    addra = 32'd36928;
    dina = {96'd0, 16'd21611, 16'd42821, 16'd59089, 16'd49166, 16'd43341, 16'd47415, 16'd45089, 16'd17852, 16'd15426, 16'd9902}; // indx = 1154
    #10;
    addra = 32'd36960;
    dina = {96'd0, 16'd55696, 16'd106, 16'd16574, 16'd3375, 16'd46267, 16'd33782, 16'd22225, 16'd29419, 16'd64974, 16'd41373}; // indx = 1155
    #10;
    addra = 32'd36992;
    dina = {96'd0, 16'd63951, 16'd21748, 16'd65433, 16'd29762, 16'd21367, 16'd23377, 16'd13721, 16'd11258, 16'd15681, 16'd33536}; // indx = 1156
    #10;
    addra = 32'd37024;
    dina = {96'd0, 16'd8185, 16'd47290, 16'd51731, 16'd16610, 16'd57718, 16'd55473, 16'd59557, 16'd10281, 16'd13149, 16'd20421}; // indx = 1157
    #10;
    addra = 32'd37056;
    dina = {96'd0, 16'd3008, 16'd52189, 16'd32920, 16'd8115, 16'd50130, 16'd41788, 16'd12529, 16'd63737, 16'd2360, 16'd55897}; // indx = 1158
    #10;
    addra = 32'd37088;
    dina = {96'd0, 16'd21620, 16'd33329, 16'd61905, 16'd63684, 16'd15466, 16'd41397, 16'd26646, 16'd58735, 16'd32573, 16'd19630}; // indx = 1159
    #10;
    addra = 32'd37120;
    dina = {96'd0, 16'd17345, 16'd27277, 16'd56486, 16'd63826, 16'd43127, 16'd23913, 16'd57912, 16'd40422, 16'd35166, 16'd6393}; // indx = 1160
    #10;
    addra = 32'd37152;
    dina = {96'd0, 16'd2408, 16'd5791, 16'd61837, 16'd1209, 16'd2966, 16'd41902, 16'd39338, 16'd23811, 16'd25982, 16'd9551}; // indx = 1161
    #10;
    addra = 32'd37184;
    dina = {96'd0, 16'd2360, 16'd61407, 16'd62783, 16'd20621, 16'd4427, 16'd36497, 16'd39335, 16'd21967, 16'd41609, 16'd6770}; // indx = 1162
    #10;
    addra = 32'd37216;
    dina = {96'd0, 16'd64982, 16'd35227, 16'd52384, 16'd54983, 16'd35475, 16'd21033, 16'd3005, 16'd59737, 16'd45939, 16'd45902}; // indx = 1163
    #10;
    addra = 32'd37248;
    dina = {96'd0, 16'd3448, 16'd12780, 16'd21462, 16'd3407, 16'd2423, 16'd9061, 16'd62844, 16'd31496, 16'd58550, 16'd54637}; // indx = 1164
    #10;
    addra = 32'd37280;
    dina = {96'd0, 16'd22554, 16'd24861, 16'd50911, 16'd17581, 16'd27183, 16'd43589, 16'd18876, 16'd33378, 16'd7002, 16'd23349}; // indx = 1165
    #10;
    addra = 32'd37312;
    dina = {96'd0, 16'd2696, 16'd61193, 16'd30182, 16'd40325, 16'd22434, 16'd46126, 16'd11312, 16'd51720, 16'd45767, 16'd35083}; // indx = 1166
    #10;
    addra = 32'd37344;
    dina = {96'd0, 16'd16900, 16'd34822, 16'd8097, 16'd10504, 16'd49617, 16'd32373, 16'd8557, 16'd52345, 16'd43907, 16'd30673}; // indx = 1167
    #10;
    addra = 32'd37376;
    dina = {96'd0, 16'd65084, 16'd11435, 16'd11513, 16'd10752, 16'd24289, 16'd23576, 16'd2267, 16'd55740, 16'd6337, 16'd22701}; // indx = 1168
    #10;
    addra = 32'd37408;
    dina = {96'd0, 16'd9748, 16'd39468, 16'd30218, 16'd45758, 16'd3510, 16'd56138, 16'd38065, 16'd31505, 16'd29664, 16'd35313}; // indx = 1169
    #10;
    addra = 32'd37440;
    dina = {96'd0, 16'd5571, 16'd31938, 16'd65047, 16'd42306, 16'd41161, 16'd40175, 16'd28277, 16'd36948, 16'd61555, 16'd50401}; // indx = 1170
    #10;
    addra = 32'd37472;
    dina = {96'd0, 16'd37480, 16'd43759, 16'd22561, 16'd8118, 16'd56237, 16'd63528, 16'd22169, 16'd19478, 16'd11103, 16'd44382}; // indx = 1171
    #10;
    addra = 32'd37504;
    dina = {96'd0, 16'd13797, 16'd11453, 16'd52363, 16'd14163, 16'd56096, 16'd64031, 16'd1225, 16'd37000, 16'd5924, 16'd17715}; // indx = 1172
    #10;
    addra = 32'd37536;
    dina = {96'd0, 16'd49681, 16'd64430, 16'd28939, 16'd58658, 16'd8662, 16'd12163, 16'd9335, 16'd63150, 16'd14998, 16'd20889}; // indx = 1173
    #10;
    addra = 32'd37568;
    dina = {96'd0, 16'd56597, 16'd20902, 16'd28882, 16'd30618, 16'd29430, 16'd15121, 16'd31828, 16'd8489, 16'd62628, 16'd3291}; // indx = 1174
    #10;
    addra = 32'd37600;
    dina = {96'd0, 16'd9306, 16'd62913, 16'd20182, 16'd44184, 16'd38126, 16'd49178, 16'd18169, 16'd54689, 16'd37156, 16'd36708}; // indx = 1175
    #10;
    addra = 32'd37632;
    dina = {96'd0, 16'd23888, 16'd54547, 16'd56214, 16'd17822, 16'd19891, 16'd54782, 16'd3924, 16'd19998, 16'd47294, 16'd41777}; // indx = 1176
    #10;
    addra = 32'd37664;
    dina = {96'd0, 16'd64066, 16'd39649, 16'd64809, 16'd46477, 16'd57210, 16'd7020, 16'd24820, 16'd58959, 16'd54141, 16'd37386}; // indx = 1177
    #10;
    addra = 32'd37696;
    dina = {96'd0, 16'd22024, 16'd15144, 16'd31872, 16'd52434, 16'd39975, 16'd8223, 16'd25448, 16'd12785, 16'd2774, 16'd19359}; // indx = 1178
    #10;
    addra = 32'd37728;
    dina = {96'd0, 16'd36447, 16'd37137, 16'd5677, 16'd43018, 16'd54122, 16'd59962, 16'd26164, 16'd52724, 16'd49020, 16'd2946}; // indx = 1179
    #10;
    addra = 32'd37760;
    dina = {96'd0, 16'd26025, 16'd50721, 16'd21202, 16'd47261, 16'd42244, 16'd10535, 16'd3811, 16'd14039, 16'd13816, 16'd41123}; // indx = 1180
    #10;
    addra = 32'd37792;
    dina = {96'd0, 16'd18614, 16'd11750, 16'd17441, 16'd16836, 16'd43959, 16'd40001, 16'd40224, 16'd5526, 16'd8912, 16'd7187}; // indx = 1181
    #10;
    addra = 32'd37824;
    dina = {96'd0, 16'd30565, 16'd33210, 16'd24823, 16'd1796, 16'd5333, 16'd2847, 16'd52271, 16'd59179, 16'd51637, 16'd11820}; // indx = 1182
    #10;
    addra = 32'd37856;
    dina = {96'd0, 16'd64473, 16'd55702, 16'd2574, 16'd33917, 16'd58385, 16'd14917, 16'd27539, 16'd25041, 16'd50870, 16'd53144}; // indx = 1183
    #10;
    addra = 32'd37888;
    dina = {96'd0, 16'd53886, 16'd27501, 16'd28336, 16'd60145, 16'd47530, 16'd3086, 16'd51241, 16'd16364, 16'd58292, 16'd63619}; // indx = 1184
    #10;
    addra = 32'd37920;
    dina = {96'd0, 16'd22880, 16'd16146, 16'd50584, 16'd16896, 16'd42983, 16'd23215, 16'd58613, 16'd39762, 16'd30327, 16'd32418}; // indx = 1185
    #10;
    addra = 32'd37952;
    dina = {96'd0, 16'd61946, 16'd22065, 16'd60599, 16'd61077, 16'd6814, 16'd18463, 16'd3450, 16'd37367, 16'd21522, 16'd38538}; // indx = 1186
    #10;
    addra = 32'd37984;
    dina = {96'd0, 16'd56126, 16'd3143, 16'd63802, 16'd47920, 16'd41692, 16'd53253, 16'd21312, 16'd36456, 16'd44496, 16'd15099}; // indx = 1187
    #10;
    addra = 32'd38016;
    dina = {96'd0, 16'd7206, 16'd19396, 16'd5679, 16'd37249, 16'd14334, 16'd54453, 16'd3201, 16'd52489, 16'd41569, 16'd34320}; // indx = 1188
    #10;
    addra = 32'd38048;
    dina = {96'd0, 16'd28259, 16'd34262, 16'd12662, 16'd18364, 16'd51543, 16'd56420, 16'd34100, 16'd56566, 16'd34279, 16'd14531}; // indx = 1189
    #10;
    addra = 32'd38080;
    dina = {96'd0, 16'd4411, 16'd65432, 16'd57413, 16'd12605, 16'd20455, 16'd22057, 16'd62292, 16'd50757, 16'd40874, 16'd28590}; // indx = 1190
    #10;
    addra = 32'd38112;
    dina = {96'd0, 16'd14933, 16'd55936, 16'd45359, 16'd24403, 16'd38294, 16'd11305, 16'd53744, 16'd56479, 16'd55680, 16'd29995}; // indx = 1191
    #10;
    addra = 32'd38144;
    dina = {96'd0, 16'd27104, 16'd62424, 16'd53594, 16'd42681, 16'd20191, 16'd38449, 16'd37430, 16'd54034, 16'd26764, 16'd901}; // indx = 1192
    #10;
    addra = 32'd38176;
    dina = {96'd0, 16'd4357, 16'd3823, 16'd32034, 16'd62980, 16'd8454, 16'd14776, 16'd41871, 16'd62206, 16'd29208, 16'd18516}; // indx = 1193
    #10;
    addra = 32'd38208;
    dina = {96'd0, 16'd54864, 16'd31628, 16'd47805, 16'd35280, 16'd56964, 16'd41734, 16'd34515, 16'd36281, 16'd42805, 16'd53271}; // indx = 1194
    #10;
    addra = 32'd38240;
    dina = {96'd0, 16'd33614, 16'd38086, 16'd51043, 16'd45544, 16'd58628, 16'd20551, 16'd50042, 16'd60145, 16'd59147, 16'd32125}; // indx = 1195
    #10;
    addra = 32'd38272;
    dina = {96'd0, 16'd38121, 16'd21904, 16'd3466, 16'd38670, 16'd1863, 16'd1877, 16'd8816, 16'd17640, 16'd28150, 16'd42108}; // indx = 1196
    #10;
    addra = 32'd38304;
    dina = {96'd0, 16'd8219, 16'd54080, 16'd14711, 16'd59847, 16'd47963, 16'd55326, 16'd20651, 16'd12007, 16'd18231, 16'd45599}; // indx = 1197
    #10;
    addra = 32'd38336;
    dina = {96'd0, 16'd54430, 16'd33003, 16'd53708, 16'd2003, 16'd55644, 16'd6362, 16'd12523, 16'd9570, 16'd35271, 16'd28752}; // indx = 1198
    #10;
    addra = 32'd38368;
    dina = {96'd0, 16'd52643, 16'd39364, 16'd32943, 16'd3584, 16'd27172, 16'd33513, 16'd33048, 16'd9344, 16'd17664, 16'd33627}; // indx = 1199
    #10;
    addra = 32'd38400;
    dina = {96'd0, 16'd53927, 16'd20569, 16'd32794, 16'd17691, 16'd32135, 16'd65463, 16'd43985, 16'd23576, 16'd60211, 16'd3233}; // indx = 1200
    #10;
    addra = 32'd38432;
    dina = {96'd0, 16'd27429, 16'd1420, 16'd50840, 16'd3595, 16'd24446, 16'd46463, 16'd23116, 16'd62581, 16'd28594, 16'd9689}; // indx = 1201
    #10;
    addra = 32'd38464;
    dina = {96'd0, 16'd63762, 16'd18220, 16'd3906, 16'd32033, 16'd49171, 16'd20030, 16'd50420, 16'd4312, 16'd54093, 16'd38503}; // indx = 1202
    #10;
    addra = 32'd38496;
    dina = {96'd0, 16'd1820, 16'd40882, 16'd15036, 16'd13338, 16'd29427, 16'd22946, 16'd56411, 16'd3239, 16'd19902, 16'd57735}; // indx = 1203
    #10;
    addra = 32'd38528;
    dina = {96'd0, 16'd633, 16'd136, 16'd3943, 16'd12786, 16'd34944, 16'd60753, 16'd61821, 16'd28760, 16'd38588, 16'd10325}; // indx = 1204
    #10;
    addra = 32'd38560;
    dina = {96'd0, 16'd28396, 16'd63380, 16'd49844, 16'd37279, 16'd60520, 16'd9766, 16'd26683, 16'd62144, 16'd34816, 16'd53922}; // indx = 1205
    #10;
    addra = 32'd38592;
    dina = {96'd0, 16'd1984, 16'd33910, 16'd42880, 16'd16611, 16'd10913, 16'd55607, 16'd22601, 16'd55525, 16'd41045, 16'd59216}; // indx = 1206
    #10;
    addra = 32'd38624;
    dina = {96'd0, 16'd39249, 16'd35786, 16'd60434, 16'd1217, 16'd48178, 16'd27090, 16'd6743, 16'd64957, 16'd31205, 16'd50931}; // indx = 1207
    #10;
    addra = 32'd38656;
    dina = {96'd0, 16'd36095, 16'd38358, 16'd33193, 16'd24728, 16'd40495, 16'd47871, 16'd18544, 16'd18661, 16'd7243, 16'd19253}; // indx = 1208
    #10;
    addra = 32'd38688;
    dina = {96'd0, 16'd64751, 16'd21555, 16'd23093, 16'd51148, 16'd32109, 16'd14190, 16'd64947, 16'd29271, 16'd63487, 16'd29056}; // indx = 1209
    #10;
    addra = 32'd38720;
    dina = {96'd0, 16'd29994, 16'd51341, 16'd43660, 16'd32140, 16'd31851, 16'd34966, 16'd4950, 16'd3801, 16'd3391, 16'd7309}; // indx = 1210
    #10;
    addra = 32'd38752;
    dina = {96'd0, 16'd33952, 16'd2615, 16'd32892, 16'd24104, 16'd18571, 16'd49932, 16'd47632, 16'd31808, 16'd53503, 16'd14224}; // indx = 1211
    #10;
    addra = 32'd38784;
    dina = {96'd0, 16'd11128, 16'd39659, 16'd37076, 16'd52984, 16'd35579, 16'd63288, 16'd1729, 16'd30778, 16'd32375, 16'd29101}; // indx = 1212
    #10;
    addra = 32'd38816;
    dina = {96'd0, 16'd33010, 16'd9106, 16'd4925, 16'd16353, 16'd4444, 16'd46085, 16'd23046, 16'd5576, 16'd42147, 16'd22676}; // indx = 1213
    #10;
    addra = 32'd38848;
    dina = {96'd0, 16'd45065, 16'd59306, 16'd16922, 16'd57524, 16'd38823, 16'd26508, 16'd26537, 16'd61725, 16'd3569, 16'd63648}; // indx = 1214
    #10;
    addra = 32'd38880;
    dina = {96'd0, 16'd205, 16'd3129, 16'd25615, 16'd36605, 16'd18315, 16'd41230, 16'd55315, 16'd26178, 16'd43165, 16'd60992}; // indx = 1215
    #10;
    addra = 32'd38912;
    dina = {96'd0, 16'd53955, 16'd10342, 16'd23172, 16'd27164, 16'd47892, 16'd29252, 16'd16996, 16'd7599, 16'd47661, 16'd34320}; // indx = 1216
    #10;
    addra = 32'd38944;
    dina = {96'd0, 16'd18525, 16'd40586, 16'd23768, 16'd31497, 16'd8424, 16'd57706, 16'd41767, 16'd52993, 16'd38443, 16'd5186}; // indx = 1217
    #10;
    addra = 32'd38976;
    dina = {96'd0, 16'd55744, 16'd60970, 16'd57668, 16'd37721, 16'd57349, 16'd24812, 16'd54221, 16'd23805, 16'd65114, 16'd18695}; // indx = 1218
    #10;
    addra = 32'd39008;
    dina = {96'd0, 16'd51726, 16'd43548, 16'd65270, 16'd13376, 16'd27992, 16'd46959, 16'd50162, 16'd27155, 16'd46391, 16'd38416}; // indx = 1219
    #10;
    addra = 32'd39040;
    dina = {96'd0, 16'd1955, 16'd48758, 16'd16275, 16'd63329, 16'd63436, 16'd39604, 16'd63786, 16'd19131, 16'd31663, 16'd63374}; // indx = 1220
    #10;
    addra = 32'd39072;
    dina = {96'd0, 16'd53805, 16'd22139, 16'd42780, 16'd20, 16'd22658, 16'd52324, 16'd39314, 16'd64676, 16'd35267, 16'd64863}; // indx = 1221
    #10;
    addra = 32'd39104;
    dina = {96'd0, 16'd17459, 16'd46198, 16'd38110, 16'd4169, 16'd28231, 16'd30375, 16'd61001, 16'd50329, 16'd20613, 16'd36072}; // indx = 1222
    #10;
    addra = 32'd39136;
    dina = {96'd0, 16'd12086, 16'd26915, 16'd3531, 16'd3181, 16'd28998, 16'd55928, 16'd17181, 16'd25175, 16'd11467, 16'd63442}; // indx = 1223
    #10;
    addra = 32'd39168;
    dina = {96'd0, 16'd60430, 16'd42301, 16'd51706, 16'd52751, 16'd59087, 16'd53881, 16'd20080, 16'd2597, 16'd19483, 16'd12271}; // indx = 1224
    #10;
    addra = 32'd39200;
    dina = {96'd0, 16'd39788, 16'd57427, 16'd44424, 16'd13299, 16'd1827, 16'd19929, 16'd40876, 16'd15030, 16'd16560, 16'd18706}; // indx = 1225
    #10;
    addra = 32'd39232;
    dina = {96'd0, 16'd39926, 16'd53255, 16'd24856, 16'd59525, 16'd27914, 16'd62098, 16'd46347, 16'd14932, 16'd8675, 16'd13850}; // indx = 1226
    #10;
    addra = 32'd39264;
    dina = {96'd0, 16'd39011, 16'd58833, 16'd17195, 16'd52101, 16'd60300, 16'd33297, 16'd28508, 16'd18875, 16'd10405, 16'd22180}; // indx = 1227
    #10;
    addra = 32'd39296;
    dina = {96'd0, 16'd31059, 16'd63627, 16'd54902, 16'd44064, 16'd31051, 16'd14733, 16'd25567, 16'd11740, 16'd61957, 16'd39859}; // indx = 1228
    #10;
    addra = 32'd39328;
    dina = {96'd0, 16'd62848, 16'd46363, 16'd16564, 16'd1129, 16'd16299, 16'd28830, 16'd53418, 16'd63349, 16'd22265, 16'd63949}; // indx = 1229
    #10;
    addra = 32'd39360;
    dina = {96'd0, 16'd41243, 16'd45587, 16'd4704, 16'd44971, 16'd44119, 16'd29024, 16'd12769, 16'd17035, 16'd2099, 16'd46940}; // indx = 1230
    #10;
    addra = 32'd39392;
    dina = {96'd0, 16'd27947, 16'd26747, 16'd29862, 16'd50314, 16'd64053, 16'd59954, 16'd15891, 16'd47050, 16'd27822, 16'd59440}; // indx = 1231
    #10;
    addra = 32'd39424;
    dina = {96'd0, 16'd21647, 16'd22312, 16'd54825, 16'd40795, 16'd11831, 16'd2110, 16'd39138, 16'd22215, 16'd15808, 16'd41546}; // indx = 1232
    #10;
    addra = 32'd39456;
    dina = {96'd0, 16'd8646, 16'd57984, 16'd5273, 16'd64054, 16'd44623, 16'd35659, 16'd30166, 16'd31870, 16'd29987, 16'd48299}; // indx = 1233
    #10;
    addra = 32'd39488;
    dina = {96'd0, 16'd18031, 16'd40563, 16'd10566, 16'd9355, 16'd43678, 16'd34157, 16'd13510, 16'd59668, 16'd56986, 16'd21390}; // indx = 1234
    #10;
    addra = 32'd39520;
    dina = {96'd0, 16'd17168, 16'd60431, 16'd6559, 16'd55971, 16'd56861, 16'd18986, 16'd13407, 16'd44163, 16'd23463, 16'd4075}; // indx = 1235
    #10;
    addra = 32'd39552;
    dina = {96'd0, 16'd5162, 16'd62902, 16'd40946, 16'd505, 16'd47788, 16'd49050, 16'd17644, 16'd38833, 16'd26651, 16'd13624}; // indx = 1236
    #10;
    addra = 32'd39584;
    dina = {96'd0, 16'd62900, 16'd33753, 16'd2958, 16'd48694, 16'd44915, 16'd25527, 16'd6961, 16'd19386, 16'd23938, 16'd57644}; // indx = 1237
    #10;
    addra = 32'd39616;
    dina = {96'd0, 16'd51643, 16'd58512, 16'd37745, 16'd25610, 16'd37280, 16'd65085, 16'd7144, 16'd62231, 16'd35975, 16'd28157}; // indx = 1238
    #10;
    addra = 32'd39648;
    dina = {96'd0, 16'd20201, 16'd8747, 16'd47112, 16'd8781, 16'd1107, 16'd62352, 16'd4534, 16'd57117, 16'd8218, 16'd32496}; // indx = 1239
    #10;
    addra = 32'd39680;
    dina = {96'd0, 16'd52060, 16'd15635, 16'd38963, 16'd56426, 16'd62773, 16'd45557, 16'd20635, 16'd31355, 16'd51622, 16'd14381}; // indx = 1240
    #10;
    addra = 32'd39712;
    dina = {96'd0, 16'd49941, 16'd3218, 16'd27400, 16'd64335, 16'd22840, 16'd32251, 16'd137, 16'd25850, 16'd62071, 16'd42188}; // indx = 1241
    #10;
    addra = 32'd39744;
    dina = {96'd0, 16'd804, 16'd20337, 16'd43392, 16'd14260, 16'd11979, 16'd23196, 16'd50396, 16'd26606, 16'd62397, 16'd39412}; // indx = 1242
    #10;
    addra = 32'd39776;
    dina = {96'd0, 16'd7907, 16'd24719, 16'd5034, 16'd9154, 16'd29649, 16'd37466, 16'd399, 16'd51335, 16'd5624, 16'd17019}; // indx = 1243
    #10;
    addra = 32'd39808;
    dina = {96'd0, 16'd4674, 16'd42745, 16'd63511, 16'd35380, 16'd10617, 16'd20333, 16'd13939, 16'd16388, 16'd21579, 16'd40015}; // indx = 1244
    #10;
    addra = 32'd39840;
    dina = {96'd0, 16'd36450, 16'd25633, 16'd9226, 16'd52314, 16'd59606, 16'd55118, 16'd54687, 16'd19257, 16'd12936, 16'd61624}; // indx = 1245
    #10;
    addra = 32'd39872;
    dina = {96'd0, 16'd39751, 16'd14016, 16'd31016, 16'd27362, 16'd32808, 16'd59905, 16'd46412, 16'd55437, 16'd44930, 16'd29154}; // indx = 1246
    #10;
    addra = 32'd39904;
    dina = {96'd0, 16'd5660, 16'd48431, 16'd32081, 16'd28573, 16'd31473, 16'd22263, 16'd52039, 16'd50373, 16'd26912, 16'd22372}; // indx = 1247
    #10;
    addra = 32'd39936;
    dina = {96'd0, 16'd19916, 16'd41726, 16'd52141, 16'd52367, 16'd43042, 16'd28542, 16'd60825, 16'd12214, 16'd48667, 16'd23315}; // indx = 1248
    #10;
    addra = 32'd39968;
    dina = {96'd0, 16'd44653, 16'd7340, 16'd19293, 16'd26996, 16'd44313, 16'd61085, 16'd1502, 16'd52147, 16'd57091, 16'd41882}; // indx = 1249
    #10;
    addra = 32'd40000;
    dina = {96'd0, 16'd19808, 16'd30757, 16'd16409, 16'd27578, 16'd6610, 16'd64182, 16'd60025, 16'd28021, 16'd50710, 16'd45644}; // indx = 1250
    #10;
    addra = 32'd40032;
    dina = {96'd0, 16'd55754, 16'd45782, 16'd36835, 16'd49714, 16'd20206, 16'd60256, 16'd31719, 16'd12281, 16'd43960, 16'd50645}; // indx = 1251
    #10;
    addra = 32'd40064;
    dina = {96'd0, 16'd50356, 16'd43651, 16'd60872, 16'd20874, 16'd45787, 16'd13568, 16'd48723, 16'd26442, 16'd55218, 16'd2468}; // indx = 1252
    #10;
    addra = 32'd40096;
    dina = {96'd0, 16'd47107, 16'd5119, 16'd4409, 16'd30794, 16'd10573, 16'd37359, 16'd64223, 16'd13892, 16'd13009, 16'd14959}; // indx = 1253
    #10;
    addra = 32'd40128;
    dina = {96'd0, 16'd7894, 16'd48193, 16'd25016, 16'd32208, 16'd55979, 16'd7731, 16'd5378, 16'd23402, 16'd3071, 16'd62185}; // indx = 1254
    #10;
    addra = 32'd40160;
    dina = {96'd0, 16'd4479, 16'd45239, 16'd45949, 16'd1036, 16'd12236, 16'd61352, 16'd54285, 16'd39457, 16'd3156, 16'd1660}; // indx = 1255
    #10;
    addra = 32'd40192;
    dina = {96'd0, 16'd1550, 16'd12474, 16'd59656, 16'd6247, 16'd22008, 16'd32008, 16'd61258, 16'd4279, 16'd46947, 16'd35789}; // indx = 1256
    #10;
    addra = 32'd40224;
    dina = {96'd0, 16'd14128, 16'd56655, 16'd39051, 16'd62309, 16'd4729, 16'd44235, 16'd7435, 16'd55275, 16'd44104, 16'd61797}; // indx = 1257
    #10;
    addra = 32'd40256;
    dina = {96'd0, 16'd7071, 16'd44170, 16'd44961, 16'd43920, 16'd4568, 16'd48828, 16'd5321, 16'd15187, 16'd52537, 16'd48137}; // indx = 1258
    #10;
    addra = 32'd40288;
    dina = {96'd0, 16'd29280, 16'd55298, 16'd20995, 16'd62040, 16'd4640, 16'd51998, 16'd21527, 16'd51420, 16'd30681, 16'd34887}; // indx = 1259
    #10;
    addra = 32'd40320;
    dina = {96'd0, 16'd53868, 16'd62789, 16'd26311, 16'd62504, 16'd57010, 16'd60851, 16'd16343, 16'd7565, 16'd57009, 16'd21810}; // indx = 1260
    #10;
    addra = 32'd40352;
    dina = {96'd0, 16'd51576, 16'd25064, 16'd19158, 16'd25401, 16'd10199, 16'd55345, 16'd2213, 16'd59819, 16'd9810, 16'd14118}; // indx = 1261
    #10;
    addra = 32'd40384;
    dina = {96'd0, 16'd19487, 16'd9304, 16'd10773, 16'd38077, 16'd33692, 16'd23011, 16'd27240, 16'd25798, 16'd7746, 16'd54363}; // indx = 1262
    #10;
    addra = 32'd40416;
    dina = {96'd0, 16'd56678, 16'd7342, 16'd37088, 16'd16049, 16'd20110, 16'd40145, 16'd13424, 16'd39134, 16'd1539, 16'd48991}; // indx = 1263
    #10;
    addra = 32'd40448;
    dina = {96'd0, 16'd3505, 16'd2741, 16'd54742, 16'd46774, 16'd41961, 16'd24236, 16'd21961, 16'd56585, 16'd16045, 16'd63198}; // indx = 1264
    #10;
    addra = 32'd40480;
    dina = {96'd0, 16'd14136, 16'd47169, 16'd5357, 16'd33567, 16'd19372, 16'd56004, 16'd17627, 16'd47279, 16'd24539, 16'd19251}; // indx = 1265
    #10;
    addra = 32'd40512;
    dina = {96'd0, 16'd34632, 16'd7225, 16'd9558, 16'd6555, 16'd58901, 16'd63388, 16'd51090, 16'd16102, 16'd60216, 16'd23288}; // indx = 1266
    #10;
    addra = 32'd40544;
    dina = {96'd0, 16'd22300, 16'd55904, 16'd39500, 16'd60825, 16'd63724, 16'd33698, 16'd20795, 16'd25790, 16'd17124, 16'd45630}; // indx = 1267
    #10;
    addra = 32'd40576;
    dina = {96'd0, 16'd12367, 16'd62348, 16'd51588, 16'd24119, 16'd42744, 16'd7076, 16'd64052, 16'd6201, 16'd51816, 16'd37935}; // indx = 1268
    #10;
    addra = 32'd40608;
    dina = {96'd0, 16'd52245, 16'd4248, 16'd48810, 16'd25757, 16'd55144, 16'd2534, 16'd57609, 16'd49838, 16'd37205, 16'd65028}; // indx = 1269
    #10;
    addra = 32'd40640;
    dina = {96'd0, 16'd59324, 16'd45441, 16'd49075, 16'd14327, 16'd56975, 16'd33257, 16'd26068, 16'd6279, 16'd15675, 16'd34027}; // indx = 1270
    #10;
    addra = 32'd40672;
    dina = {96'd0, 16'd31667, 16'd576, 16'd5080, 16'd57637, 16'd11125, 16'd7743, 16'd30643, 16'd24227, 16'd22229, 16'd19108}; // indx = 1271
    #10;
    addra = 32'd40704;
    dina = {96'd0, 16'd46126, 16'd28887, 16'd56968, 16'd49395, 16'd14780, 16'd49143, 16'd51528, 16'd63365, 16'd5025, 16'd2795}; // indx = 1272
    #10;
    addra = 32'd40736;
    dina = {96'd0, 16'd55384, 16'd27239, 16'd35235, 16'd26533, 16'd34231, 16'd4334, 16'd49949, 16'd52019, 16'd25415, 16'd48190}; // indx = 1273
    #10;
    addra = 32'd40768;
    dina = {96'd0, 16'd48198, 16'd6482, 16'd52020, 16'd11524, 16'd20547, 16'd48720, 16'd46219, 16'd51069, 16'd8959, 16'd56960}; // indx = 1274
    #10;
    addra = 32'd40800;
    dina = {96'd0, 16'd30405, 16'd15981, 16'd6807, 16'd8624, 16'd23442, 16'd58176, 16'd50765, 16'd30001, 16'd51749, 16'd58709}; // indx = 1275
    #10;
    addra = 32'd40832;
    dina = {96'd0, 16'd12202, 16'd24116, 16'd30609, 16'd31973, 16'd54189, 16'd38275, 16'd14218, 16'd39654, 16'd60041, 16'd21725}; // indx = 1276
    #10;
    addra = 32'd40864;
    dina = {96'd0, 16'd12315, 16'd31368, 16'd863, 16'd35529, 16'd55444, 16'd40484, 16'd38523, 16'd15243, 16'd41103, 16'd47703}; // indx = 1277
    #10;
    addra = 32'd40896;
    dina = {96'd0, 16'd4967, 16'd51988, 16'd17076, 16'd48664, 16'd31110, 16'd9411, 16'd2185, 16'd47128, 16'd22126, 16'd33031}; // indx = 1278
    #10;
    addra = 32'd40928;
    dina = {96'd0, 16'd62036, 16'd46249, 16'd5686, 16'd57434, 16'd42334, 16'd7920, 16'd20103, 16'd55298, 16'd49870, 16'd54456}; // indx = 1279
    #10;
    addra = 32'd40960;
    dina = {96'd0, 16'd29799, 16'd35355, 16'd28942, 16'd20859, 16'd39750, 16'd34173, 16'd8419, 16'd40141, 16'd904, 16'd8018}; // indx = 1280
    #10;
    addra = 32'd40992;
    dina = {96'd0, 16'd64130, 16'd32440, 16'd2443, 16'd25817, 16'd9247, 16'd41068, 16'd39543, 16'd25662, 16'd33029, 16'd1398}; // indx = 1281
    #10;
    addra = 32'd41024;
    dina = {96'd0, 16'd65171, 16'd58627, 16'd13398, 16'd9678, 16'd29807, 16'd57616, 16'd11527, 16'd36690, 16'd20177, 16'd58606}; // indx = 1282
    #10;
    addra = 32'd41056;
    dina = {96'd0, 16'd54783, 16'd29227, 16'd60704, 16'd63380, 16'd22775, 16'd61146, 16'd58509, 16'd39607, 16'd43328, 16'd6682}; // indx = 1283
    #10;
    addra = 32'd41088;
    dina = {96'd0, 16'd37428, 16'd44645, 16'd3829, 16'd64177, 16'd12919, 16'd47718, 16'd50330, 16'd7768, 16'd53326, 16'd37383}; // indx = 1284
    #10;
    addra = 32'd41120;
    dina = {96'd0, 16'd61578, 16'd50486, 16'd5047, 16'd12286, 16'd47125, 16'd47551, 16'd49389, 16'd10691, 16'd46390, 16'd157}; // indx = 1285
    #10;
    addra = 32'd41152;
    dina = {96'd0, 16'd9139, 16'd59654, 16'd54387, 16'd24627, 16'd14166, 16'd30526, 16'd42137, 16'd26297, 16'd50974, 16'd45828}; // indx = 1286
    #10;
    addra = 32'd41184;
    dina = {96'd0, 16'd2554, 16'd32747, 16'd9811, 16'd45840, 16'd35789, 16'd19746, 16'd49026, 16'd43502, 16'd8603, 16'd37952}; // indx = 1287
    #10;
    addra = 32'd41216;
    dina = {96'd0, 16'd17927, 16'd13892, 16'd54907, 16'd20126, 16'd53817, 16'd2763, 16'd64077, 16'd43794, 16'd61687, 16'd50611}; // indx = 1288
    #10;
    addra = 32'd41248;
    dina = {96'd0, 16'd48060, 16'd6366, 16'd48209, 16'd19667, 16'd20839, 16'd52001, 16'd23477, 16'd49193, 16'd9280, 16'd40114}; // indx = 1289
    #10;
    addra = 32'd41280;
    dina = {96'd0, 16'd42814, 16'd11475, 16'd23647, 16'd22668, 16'd23808, 16'd53381, 16'd39816, 16'd61403, 16'd10035, 16'd40634}; // indx = 1290
    #10;
    addra = 32'd41312;
    dina = {96'd0, 16'd38417, 16'd4939, 16'd39564, 16'd40610, 16'd1107, 16'd28549, 16'd30428, 16'd25643, 16'd50597, 16'd26622}; // indx = 1291
    #10;
    addra = 32'd41344;
    dina = {96'd0, 16'd45263, 16'd38147, 16'd16399, 16'd37948, 16'd4858, 16'd32237, 16'd9041, 16'd37045, 16'd1154, 16'd30217}; // indx = 1292
    #10;
    addra = 32'd41376;
    dina = {96'd0, 16'd60534, 16'd42201, 16'd37084, 16'd27490, 16'd1628, 16'd25505, 16'd12237, 16'd18029, 16'd30236, 16'd1742}; // indx = 1293
    #10;
    addra = 32'd41408;
    dina = {96'd0, 16'd17121, 16'd11503, 16'd47779, 16'd19141, 16'd10289, 16'd46507, 16'd15849, 16'd24827, 16'd60471, 16'd43637}; // indx = 1294
    #10;
    addra = 32'd41440;
    dina = {96'd0, 16'd14503, 16'd22576, 16'd15627, 16'd33919, 16'd63978, 16'd64876, 16'd47563, 16'd4678, 16'd2439, 16'd18460}; // indx = 1295
    #10;
    addra = 32'd41472;
    dina = {96'd0, 16'd34374, 16'd551, 16'd59529, 16'd36076, 16'd58485, 16'd36378, 16'd25668, 16'd51272, 16'd47643, 16'd16572}; // indx = 1296
    #10;
    addra = 32'd41504;
    dina = {96'd0, 16'd55318, 16'd39090, 16'd19510, 16'd41436, 16'd38786, 16'd51816, 16'd5084, 16'd795, 16'd61032, 16'd64407}; // indx = 1297
    #10;
    addra = 32'd41536;
    dina = {96'd0, 16'd58484, 16'd61284, 16'd56160, 16'd62400, 16'd16032, 16'd43034, 16'd51850, 16'd43686, 16'd50921, 16'd59421}; // indx = 1298
    #10;
    addra = 32'd41568;
    dina = {96'd0, 16'd32808, 16'd10574, 16'd52336, 16'd23471, 16'd6133, 16'd49638, 16'd55627, 16'd12031, 16'd8522, 16'd35219}; // indx = 1299
    #10;
    addra = 32'd41600;
    dina = {96'd0, 16'd60633, 16'd45779, 16'd60610, 16'd16065, 16'd2260, 16'd34575, 16'd5391, 16'd57016, 16'd34983, 16'd54139}; // indx = 1300
    #10;
    addra = 32'd41632;
    dina = {96'd0, 16'd20683, 16'd34603, 16'd8650, 16'd41188, 16'd22226, 16'd1401, 16'd3849, 16'd20770, 16'd35808, 16'd45219}; // indx = 1301
    #10;
    addra = 32'd41664;
    dina = {96'd0, 16'd40564, 16'd55433, 16'd33247, 16'd25834, 16'd48018, 16'd48621, 16'd45772, 16'd24425, 16'd18435, 16'd7747}; // indx = 1302
    #10;
    addra = 32'd41696;
    dina = {96'd0, 16'd53604, 16'd10211, 16'd34186, 16'd47429, 16'd19724, 16'd14789, 16'd30670, 16'd52636, 16'd12135, 16'd2970}; // indx = 1303
    #10;
    addra = 32'd41728;
    dina = {96'd0, 16'd65100, 16'd50667, 16'd40604, 16'd38560, 16'd54378, 16'd29440, 16'd25911, 16'd35792, 16'd27456, 16'd25563}; // indx = 1304
    #10;
    addra = 32'd41760;
    dina = {96'd0, 16'd55557, 16'd5757, 16'd60326, 16'd18299, 16'd60246, 16'd20894, 16'd35055, 16'd44438, 16'd51342, 16'd15632}; // indx = 1305
    #10;
    addra = 32'd41792;
    dina = {96'd0, 16'd19710, 16'd23047, 16'd35773, 16'd24268, 16'd17761, 16'd20756, 16'd16902, 16'd5261, 16'd5249, 16'd43267}; // indx = 1306
    #10;
    addra = 32'd41824;
    dina = {96'd0, 16'd54351, 16'd41746, 16'd5376, 16'd8243, 16'd32686, 16'd59405, 16'd29182, 16'd61827, 16'd3541, 16'd41735}; // indx = 1307
    #10;
    addra = 32'd41856;
    dina = {96'd0, 16'd15703, 16'd38954, 16'd46663, 16'd35500, 16'd12817, 16'd61231, 16'd20968, 16'd40853, 16'd41452, 16'd59112}; // indx = 1308
    #10;
    addra = 32'd41888;
    dina = {96'd0, 16'd5059, 16'd58618, 16'd49337, 16'd41293, 16'd41362, 16'd6048, 16'd28589, 16'd4728, 16'd1593, 16'd63923}; // indx = 1309
    #10;
    addra = 32'd41920;
    dina = {96'd0, 16'd28518, 16'd38536, 16'd26088, 16'd38513, 16'd11865, 16'd18758, 16'd48253, 16'd43798, 16'd25499, 16'd10946}; // indx = 1310
    #10;
    addra = 32'd41952;
    dina = {96'd0, 16'd25838, 16'd36161, 16'd64969, 16'd32546, 16'd43127, 16'd27801, 16'd26397, 16'd7181, 16'd22480, 16'd3510}; // indx = 1311
    #10;
    addra = 32'd41984;
    dina = {96'd0, 16'd45008, 16'd13640, 16'd24240, 16'd25809, 16'd23943, 16'd62816, 16'd64516, 16'd55920, 16'd46777, 16'd58711}; // indx = 1312
    #10;
    addra = 32'd42016;
    dina = {96'd0, 16'd10967, 16'd21249, 16'd50768, 16'd27323, 16'd9244, 16'd61816, 16'd29302, 16'd47076, 16'd48642, 16'd18715}; // indx = 1313
    #10;
    addra = 32'd42048;
    dina = {96'd0, 16'd127, 16'd25837, 16'd29141, 16'd5774, 16'd18868, 16'd23583, 16'd697, 16'd20087, 16'd24226, 16'd61107}; // indx = 1314
    #10;
    addra = 32'd42080;
    dina = {96'd0, 16'd4840, 16'd3330, 16'd31512, 16'd25041, 16'd22535, 16'd8702, 16'd51917, 16'd51786, 16'd45146, 16'd35641}; // indx = 1315
    #10;
    addra = 32'd42112;
    dina = {96'd0, 16'd23991, 16'd49296, 16'd43855, 16'd42365, 16'd58778, 16'd41207, 16'd51108, 16'd1239, 16'd35484, 16'd63659}; // indx = 1316
    #10;
    addra = 32'd42144;
    dina = {96'd0, 16'd36248, 16'd29200, 16'd52257, 16'd9225, 16'd40051, 16'd50705, 16'd8565, 16'd6388, 16'd39764, 16'd26325}; // indx = 1317
    #10;
    addra = 32'd42176;
    dina = {96'd0, 16'd38178, 16'd36498, 16'd55414, 16'd44151, 16'd3838, 16'd39635, 16'd5967, 16'd10468, 16'd3917, 16'd36404}; // indx = 1318
    #10;
    addra = 32'd42208;
    dina = {96'd0, 16'd28676, 16'd21509, 16'd45029, 16'd55400, 16'd44872, 16'd32694, 16'd6053, 16'd59216, 16'd51411, 16'd41650}; // indx = 1319
    #10;
    addra = 32'd42240;
    dina = {96'd0, 16'd22811, 16'd24864, 16'd61483, 16'd30430, 16'd8450, 16'd10834, 16'd41001, 16'd31543, 16'd50894, 16'd5620}; // indx = 1320
    #10;
    addra = 32'd42272;
    dina = {96'd0, 16'd8618, 16'd36033, 16'd57458, 16'd2156, 16'd31978, 16'd62465, 16'd2189, 16'd18267, 16'd25062, 16'd54128}; // indx = 1321
    #10;
    addra = 32'd42304;
    dina = {96'd0, 16'd65501, 16'd64853, 16'd44754, 16'd57932, 16'd54688, 16'd1092, 16'd15061, 16'd60870, 16'd48640, 16'd41645}; // indx = 1322
    #10;
    addra = 32'd42336;
    dina = {96'd0, 16'd37113, 16'd305, 16'd56258, 16'd55021, 16'd41061, 16'd27730, 16'd41955, 16'd20095, 16'd62331, 16'd28902}; // indx = 1323
    #10;
    addra = 32'd42368;
    dina = {96'd0, 16'd63726, 16'd6061, 16'd47339, 16'd62200, 16'd195, 16'd45090, 16'd22045, 16'd46465, 16'd60925, 16'd43246}; // indx = 1324
    #10;
    addra = 32'd42400;
    dina = {96'd0, 16'd59844, 16'd24098, 16'd8333, 16'd61495, 16'd2553, 16'd49799, 16'd35161, 16'd16301, 16'd871, 16'd42096}; // indx = 1325
    #10;
    addra = 32'd42432;
    dina = {96'd0, 16'd35855, 16'd15836, 16'd15601, 16'd38188, 16'd39887, 16'd31789, 16'd18844, 16'd43549, 16'd15851, 16'd39962}; // indx = 1326
    #10;
    addra = 32'd42464;
    dina = {96'd0, 16'd15182, 16'd34333, 16'd42303, 16'd277, 16'd59678, 16'd5039, 16'd18932, 16'd64592, 16'd3203, 16'd19802}; // indx = 1327
    #10;
    addra = 32'd42496;
    dina = {96'd0, 16'd46954, 16'd41612, 16'd24093, 16'd46499, 16'd44967, 16'd58438, 16'd15755, 16'd24494, 16'd29284, 16'd18717}; // indx = 1328
    #10;
    addra = 32'd42528;
    dina = {96'd0, 16'd14949, 16'd39456, 16'd10175, 16'd60267, 16'd61737, 16'd28248, 16'd14654, 16'd48262, 16'd52005, 16'd39016}; // indx = 1329
    #10;
    addra = 32'd42560;
    dina = {96'd0, 16'd49237, 16'd52276, 16'd33574, 16'd11805, 16'd50293, 16'd47752, 16'd25058, 16'd62213, 16'd461, 16'd29650}; // indx = 1330
    #10;
    addra = 32'd42592;
    dina = {96'd0, 16'd57268, 16'd59527, 16'd34382, 16'd322, 16'd27634, 16'd55241, 16'd23298, 16'd55209, 16'd29361, 16'd51751}; // indx = 1331
    #10;
    addra = 32'd42624;
    dina = {96'd0, 16'd22887, 16'd4595, 16'd39215, 16'd8557, 16'd27425, 16'd15042, 16'd59036, 16'd2534, 16'd45038, 16'd21108}; // indx = 1332
    #10;
    addra = 32'd42656;
    dina = {96'd0, 16'd34186, 16'd13077, 16'd7808, 16'd41642, 16'd38712, 16'd15, 16'd46718, 16'd4584, 16'd40932, 16'd64653}; // indx = 1333
    #10;
    addra = 32'd42688;
    dina = {96'd0, 16'd50072, 16'd23679, 16'd57417, 16'd22111, 16'd20381, 16'd46779, 16'd8069, 16'd30822, 16'd23777, 16'd52919}; // indx = 1334
    #10;
    addra = 32'd42720;
    dina = {96'd0, 16'd47159, 16'd49644, 16'd23076, 16'd13073, 16'd55179, 16'd2739, 16'd32221, 16'd27699, 16'd612, 16'd29865}; // indx = 1335
    #10;
    addra = 32'd42752;
    dina = {96'd0, 16'd10006, 16'd57559, 16'd10031, 16'd42281, 16'd33972, 16'd18902, 16'd14322, 16'd24809, 16'd38575, 16'd42832}; // indx = 1336
    #10;
    addra = 32'd42784;
    dina = {96'd0, 16'd23323, 16'd48902, 16'd53575, 16'd56162, 16'd31962, 16'd17434, 16'd21614, 16'd47769, 16'd31204, 16'd41034}; // indx = 1337
    #10;
    addra = 32'd42816;
    dina = {96'd0, 16'd51653, 16'd33086, 16'd19994, 16'd62283, 16'd47912, 16'd5198, 16'd37547, 16'd31102, 16'd48251, 16'd16749}; // indx = 1338
    #10;
    addra = 32'd42848;
    dina = {96'd0, 16'd3615, 16'd21238, 16'd35748, 16'd1041, 16'd27172, 16'd11416, 16'd56963, 16'd28514, 16'd63142, 16'd35810}; // indx = 1339
    #10;
    addra = 32'd42880;
    dina = {96'd0, 16'd50828, 16'd52546, 16'd65279, 16'd60744, 16'd57023, 16'd56676, 16'd59277, 16'd7331, 16'd30053, 16'd44411}; // indx = 1340
    #10;
    addra = 32'd42912;
    dina = {96'd0, 16'd8169, 16'd24704, 16'd60354, 16'd24542, 16'd7663, 16'd37815, 16'd47214, 16'd20512, 16'd43250, 16'd28269}; // indx = 1341
    #10;
    addra = 32'd42944;
    dina = {96'd0, 16'd17035, 16'd6392, 16'd60885, 16'd17924, 16'd53644, 16'd4677, 16'd62960, 16'd50047, 16'd3212, 16'd63646}; // indx = 1342
    #10;
    addra = 32'd42976;
    dina = {96'd0, 16'd10450, 16'd31095, 16'd59907, 16'd42404, 16'd1298, 16'd33189, 16'd60044, 16'd62100, 16'd8764, 16'd49934}; // indx = 1343
    #10;
    addra = 32'd43008;
    dina = {96'd0, 16'd47709, 16'd60333, 16'd55711, 16'd26199, 16'd55568, 16'd57250, 16'd1491, 16'd35497, 16'd47198, 16'd34124}; // indx = 1344
    #10;
    addra = 32'd43040;
    dina = {96'd0, 16'd24714, 16'd19410, 16'd8700, 16'd35940, 16'd19727, 16'd40640, 16'd49657, 16'd26306, 16'd58572, 16'd61930}; // indx = 1345
    #10;
    addra = 32'd43072;
    dina = {96'd0, 16'd63544, 16'd45355, 16'd17054, 16'd47256, 16'd4606, 16'd14552, 16'd39099, 16'd1062, 16'd18297, 16'd52055}; // indx = 1346
    #10;
    addra = 32'd43104;
    dina = {96'd0, 16'd32751, 16'd38395, 16'd9651, 16'd39314, 16'd27199, 16'd7556, 16'd27667, 16'd55963, 16'd13482, 16'd35412}; // indx = 1347
    #10;
    addra = 32'd43136;
    dina = {96'd0, 16'd31372, 16'd63970, 16'd497, 16'd59519, 16'd58674, 16'd25972, 16'd35441, 16'd12695, 16'd15656, 16'd28254}; // indx = 1348
    #10;
    addra = 32'd43168;
    dina = {96'd0, 16'd64295, 16'd14813, 16'd42515, 16'd46981, 16'd5173, 16'd50914, 16'd34419, 16'd56540, 16'd49123, 16'd57171}; // indx = 1349
    #10;
    addra = 32'd43200;
    dina = {96'd0, 16'd23105, 16'd6248, 16'd30268, 16'd41425, 16'd62551, 16'd18663, 16'd32483, 16'd23966, 16'd9101, 16'd52594}; // indx = 1350
    #10;
    addra = 32'd43232;
    dina = {96'd0, 16'd36533, 16'd6067, 16'd28709, 16'd16830, 16'd22017, 16'd29276, 16'd35966, 16'd25517, 16'd6609, 16'd3901}; // indx = 1351
    #10;
    addra = 32'd43264;
    dina = {96'd0, 16'd40045, 16'd64876, 16'd44858, 16'd46048, 16'd1895, 16'd56405, 16'd23155, 16'd6905, 16'd19890, 16'd1860}; // indx = 1352
    #10;
    addra = 32'd43296;
    dina = {96'd0, 16'd23237, 16'd19614, 16'd8253, 16'd2706, 16'd44532, 16'd58612, 16'd28261, 16'd13884, 16'd58163, 16'd29115}; // indx = 1353
    #10;
    addra = 32'd43328;
    dina = {96'd0, 16'd4303, 16'd38939, 16'd3428, 16'd51636, 16'd58758, 16'd21668, 16'd40195, 16'd51284, 16'd39469, 16'd13459}; // indx = 1354
    #10;
    addra = 32'd43360;
    dina = {96'd0, 16'd25571, 16'd52260, 16'd20685, 16'd6187, 16'd52033, 16'd14032, 16'd47140, 16'd28253, 16'd21321, 16'd41327}; // indx = 1355
    #10;
    addra = 32'd43392;
    dina = {96'd0, 16'd50345, 16'd64884, 16'd6489, 16'd30812, 16'd18723, 16'd12, 16'd58324, 16'd45937, 16'd20017, 16'd53540}; // indx = 1356
    #10;
    addra = 32'd43424;
    dina = {96'd0, 16'd12904, 16'd44766, 16'd52345, 16'd38015, 16'd50258, 16'd22939, 16'd52269, 16'd26010, 16'd43856, 16'd26772}; // indx = 1357
    #10;
    addra = 32'd43456;
    dina = {96'd0, 16'd33032, 16'd24180, 16'd46896, 16'd4352, 16'd5846, 16'd56650, 16'd46658, 16'd24891, 16'd50958, 16'd41065}; // indx = 1358
    #10;
    addra = 32'd43488;
    dina = {96'd0, 16'd64647, 16'd28495, 16'd21606, 16'd46180, 16'd56393, 16'd61992, 16'd810, 16'd58209, 16'd27010, 16'd63429}; // indx = 1359
    #10;
    addra = 32'd43520;
    dina = {96'd0, 16'd49537, 16'd41490, 16'd39964, 16'd18375, 16'd6814, 16'd59615, 16'd61401, 16'd42669, 16'd15627, 16'd18462}; // indx = 1360
    #10;
    addra = 32'd43552;
    dina = {96'd0, 16'd8747, 16'd44669, 16'd3371, 16'd15011, 16'd53722, 16'd57618, 16'd56215, 16'd20184, 16'd47648, 16'd4863}; // indx = 1361
    #10;
    addra = 32'd43584;
    dina = {96'd0, 16'd52890, 16'd14428, 16'd37498, 16'd49628, 16'd12898, 16'd18783, 16'd19258, 16'd59141, 16'd56665, 16'd3642}; // indx = 1362
    #10;
    addra = 32'd43616;
    dina = {96'd0, 16'd52018, 16'd52828, 16'd42592, 16'd13164, 16'd56437, 16'd9020, 16'd16357, 16'd1578, 16'd51284, 16'd5793}; // indx = 1363
    #10;
    addra = 32'd43648;
    dina = {96'd0, 16'd48602, 16'd43517, 16'd5924, 16'd47229, 16'd53865, 16'd18350, 16'd32531, 16'd54708, 16'd36463, 16'd34395}; // indx = 1364
    #10;
    addra = 32'd43680;
    dina = {96'd0, 16'd30701, 16'd50527, 16'd51796, 16'd56078, 16'd36069, 16'd37134, 16'd4096, 16'd23083, 16'd14351, 16'd41774}; // indx = 1365
    #10;
    addra = 32'd43712;
    dina = {96'd0, 16'd16299, 16'd35576, 16'd3614, 16'd27571, 16'd4481, 16'd56355, 16'd11586, 16'd10046, 16'd6630, 16'd5101}; // indx = 1366
    #10;
    addra = 32'd43744;
    dina = {96'd0, 16'd51323, 16'd17848, 16'd3222, 16'd30699, 16'd30589, 16'd13133, 16'd3307, 16'd8983, 16'd38511, 16'd34084}; // indx = 1367
    #10;
    addra = 32'd43776;
    dina = {96'd0, 16'd32074, 16'd34981, 16'd8081, 16'd51888, 16'd27922, 16'd57167, 16'd52614, 16'd23095, 16'd15761, 16'd13453}; // indx = 1368
    #10;
    addra = 32'd43808;
    dina = {96'd0, 16'd2451, 16'd5970, 16'd13235, 16'd11080, 16'd28339, 16'd10413, 16'd52089, 16'd28732, 16'd31971, 16'd1268}; // indx = 1369
    #10;
    addra = 32'd43840;
    dina = {96'd0, 16'd23160, 16'd3122, 16'd62171, 16'd32872, 16'd36648, 16'd57875, 16'd377, 16'd46342, 16'd17494, 16'd58420}; // indx = 1370
    #10;
    addra = 32'd43872;
    dina = {96'd0, 16'd46218, 16'd17581, 16'd42416, 16'd13679, 16'd3425, 16'd49310, 16'd37354, 16'd48432, 16'd31966, 16'd43033}; // indx = 1371
    #10;
    addra = 32'd43904;
    dina = {96'd0, 16'd2265, 16'd54585, 16'd3976, 16'd35186, 16'd11757, 16'd36034, 16'd51409, 16'd4439, 16'd52297, 16'd13049}; // indx = 1372
    #10;
    addra = 32'd43936;
    dina = {96'd0, 16'd35305, 16'd10260, 16'd56112, 16'd2681, 16'd48758, 16'd47065, 16'd32537, 16'd46396, 16'd58075, 16'd48999}; // indx = 1373
    #10;
    addra = 32'd43968;
    dina = {96'd0, 16'd65386, 16'd18726, 16'd43121, 16'd15884, 16'd2223, 16'd34245, 16'd6930, 16'd8576, 16'd61022, 16'd60308}; // indx = 1374
    #10;
    addra = 32'd44000;
    dina = {96'd0, 16'd63674, 16'd54092, 16'd7923, 16'd26692, 16'd36015, 16'd53960, 16'd8220, 16'd31318, 16'd4022, 16'd61257}; // indx = 1375
    #10;
    addra = 32'd44032;
    dina = {96'd0, 16'd62516, 16'd24869, 16'd52698, 16'd46845, 16'd10693, 16'd12225, 16'd47037, 16'd45691, 16'd6561, 16'd17486}; // indx = 1376
    #10;
    addra = 32'd44064;
    dina = {96'd0, 16'd13580, 16'd63606, 16'd12640, 16'd6353, 16'd36746, 16'd61035, 16'd28122, 16'd13067, 16'd24242, 16'd14768}; // indx = 1377
    #10;
    addra = 32'd44096;
    dina = {96'd0, 16'd12, 16'd6835, 16'd18837, 16'd54499, 16'd26156, 16'd47271, 16'd24108, 16'd28525, 16'd19630, 16'd63260}; // indx = 1378
    #10;
    addra = 32'd44128;
    dina = {96'd0, 16'd20098, 16'd40196, 16'd27308, 16'd321, 16'd46146, 16'd54654, 16'd37105, 16'd57255, 16'd19809, 16'd222}; // indx = 1379
    #10;
    addra = 32'd44160;
    dina = {96'd0, 16'd25022, 16'd37914, 16'd31412, 16'd41213, 16'd46080, 16'd21693, 16'd12514, 16'd49487, 16'd34072, 16'd4257}; // indx = 1380
    #10;
    addra = 32'd44192;
    dina = {96'd0, 16'd19854, 16'd17032, 16'd21346, 16'd7322, 16'd28962, 16'd2475, 16'd1589, 16'd63518, 16'd499, 16'd29007}; // indx = 1381
    #10;
    addra = 32'd44224;
    dina = {96'd0, 16'd4157, 16'd1953, 16'd16700, 16'd35419, 16'd27532, 16'd38928, 16'd53836, 16'd62397, 16'd12217, 16'd8334}; // indx = 1382
    #10;
    addra = 32'd44256;
    dina = {96'd0, 16'd46771, 16'd39089, 16'd55825, 16'd53725, 16'd38558, 16'd11514, 16'd48613, 16'd41128, 16'd55663, 16'd41117}; // indx = 1383
    #10;
    addra = 32'd44288;
    dina = {96'd0, 16'd4826, 16'd36915, 16'd28715, 16'd9863, 16'd36264, 16'd3541, 16'd11932, 16'd45072, 16'd40855, 16'd58489}; // indx = 1384
    #10;
    addra = 32'd44320;
    dina = {96'd0, 16'd1774, 16'd2427, 16'd54286, 16'd55418, 16'd34079, 16'd10813, 16'd45438, 16'd37460, 16'd57380, 16'd6221}; // indx = 1385
    #10;
    addra = 32'd44352;
    dina = {96'd0, 16'd32216, 16'd60700, 16'd57840, 16'd3041, 16'd31649, 16'd3083, 16'd33558, 16'd10119, 16'd44203, 16'd46911}; // indx = 1386
    #10;
    addra = 32'd44384;
    dina = {96'd0, 16'd20474, 16'd37667, 16'd53367, 16'd11289, 16'd18949, 16'd28027, 16'd11459, 16'd4762, 16'd33433, 16'd61575}; // indx = 1387
    #10;
    addra = 32'd44416;
    dina = {96'd0, 16'd57992, 16'd35127, 16'd9786, 16'd38331, 16'd45483, 16'd25057, 16'd64285, 16'd2646, 16'd51014, 16'd6099}; // indx = 1388
    #10;
    addra = 32'd44448;
    dina = {96'd0, 16'd6780, 16'd4111, 16'd9830, 16'd32650, 16'd132, 16'd62921, 16'd10904, 16'd16145, 16'd32128, 16'd46391}; // indx = 1389
    #10;
    addra = 32'd44480;
    dina = {96'd0, 16'd1905, 16'd22531, 16'd42452, 16'd24357, 16'd26684, 16'd65148, 16'd16208, 16'd7829, 16'd2116, 16'd15466}; // indx = 1390
    #10;
    addra = 32'd44512;
    dina = {96'd0, 16'd36264, 16'd52732, 16'd64448, 16'd23014, 16'd6001, 16'd63360, 16'd7472, 16'd57645, 16'd40724, 16'd3109}; // indx = 1391
    #10;
    addra = 32'd44544;
    dina = {96'd0, 16'd32369, 16'd54542, 16'd41157, 16'd41163, 16'd49352, 16'd12956, 16'd28413, 16'd39051, 16'd20500, 16'd61922}; // indx = 1392
    #10;
    addra = 32'd44576;
    dina = {96'd0, 16'd11013, 16'd52402, 16'd33917, 16'd43142, 16'd53888, 16'd27638, 16'd31918, 16'd16376, 16'd54219, 16'd56604}; // indx = 1393
    #10;
    addra = 32'd44608;
    dina = {96'd0, 16'd29457, 16'd23062, 16'd21397, 16'd36486, 16'd24969, 16'd13419, 16'd11366, 16'd1355, 16'd13173, 16'd29743}; // indx = 1394
    #10;
    addra = 32'd44640;
    dina = {96'd0, 16'd19076, 16'd48511, 16'd28845, 16'd32741, 16'd10215, 16'd30921, 16'd64433, 16'd31883, 16'd48397, 16'd13711}; // indx = 1395
    #10;
    addra = 32'd44672;
    dina = {96'd0, 16'd39935, 16'd54797, 16'd8690, 16'd42005, 16'd41353, 16'd45224, 16'd52984, 16'd21836, 16'd30793, 16'd10312}; // indx = 1396
    #10;
    addra = 32'd44704;
    dina = {96'd0, 16'd41525, 16'd43245, 16'd5009, 16'd518, 16'd52842, 16'd32243, 16'd55012, 16'd4684, 16'd55550, 16'd46445}; // indx = 1397
    #10;
    addra = 32'd44736;
    dina = {96'd0, 16'd22911, 16'd36827, 16'd34389, 16'd20219, 16'd3227, 16'd47394, 16'd9339, 16'd7595, 16'd18270, 16'd7836}; // indx = 1398
    #10;
    addra = 32'd44768;
    dina = {96'd0, 16'd52102, 16'd14686, 16'd2000, 16'd23212, 16'd2627, 16'd44816, 16'd41054, 16'd40631, 16'd14834, 16'd39609}; // indx = 1399
    #10;
    addra = 32'd44800;
    dina = {96'd0, 16'd22661, 16'd8389, 16'd39057, 16'd53943, 16'd61132, 16'd51833, 16'd58973, 16'd17908, 16'd12612, 16'd9449}; // indx = 1400
    #10;
    addra = 32'd44832;
    dina = {96'd0, 16'd12694, 16'd15156, 16'd42117, 16'd58643, 16'd64638, 16'd12097, 16'd45417, 16'd4798, 16'd54403, 16'd42789}; // indx = 1401
    #10;
    addra = 32'd44864;
    dina = {96'd0, 16'd16144, 16'd44660, 16'd40929, 16'd17794, 16'd39464, 16'd57612, 16'd58714, 16'd31794, 16'd8765, 16'd31213}; // indx = 1402
    #10;
    addra = 32'd44896;
    dina = {96'd0, 16'd24843, 16'd2187, 16'd55191, 16'd27453, 16'd9796, 16'd32026, 16'd7690, 16'd44807, 16'd46241, 16'd64236}; // indx = 1403
    #10;
    addra = 32'd44928;
    dina = {96'd0, 16'd7653, 16'd157, 16'd52163, 16'd16299, 16'd1174, 16'd48178, 16'd44526, 16'd6685, 16'd62531, 16'd18185}; // indx = 1404
    #10;
    addra = 32'd44960;
    dina = {96'd0, 16'd41459, 16'd17314, 16'd14521, 16'd11623, 16'd7451, 16'd15910, 16'd7854, 16'd43166, 16'd62518, 16'd43327}; // indx = 1405
    #10;
    addra = 32'd44992;
    dina = {96'd0, 16'd20869, 16'd54433, 16'd24749, 16'd62042, 16'd15789, 16'd58721, 16'd6174, 16'd45068, 16'd53846, 16'd23802}; // indx = 1406
    #10;
    addra = 32'd45024;
    dina = {96'd0, 16'd3831, 16'd43625, 16'd1812, 16'd16331, 16'd40918, 16'd59453, 16'd11676, 16'd9365, 16'd54627, 16'd34036}; // indx = 1407
    #10;
    addra = 32'd45056;
    dina = {96'd0, 16'd1243, 16'd34071, 16'd43225, 16'd1717, 16'd28912, 16'd44560, 16'd17202, 16'd10809, 16'd56198, 16'd19678}; // indx = 1408
    #10;
    addra = 32'd45088;
    dina = {96'd0, 16'd63444, 16'd31915, 16'd62306, 16'd61768, 16'd22968, 16'd34809, 16'd48831, 16'd30157, 16'd25281, 16'd50359}; // indx = 1409
    #10;
    addra = 32'd45120;
    dina = {96'd0, 16'd13648, 16'd44264, 16'd36291, 16'd31209, 16'd22061, 16'd48929, 16'd56616, 16'd554, 16'd23361, 16'd25013}; // indx = 1410
    #10;
    addra = 32'd45152;
    dina = {96'd0, 16'd1248, 16'd10612, 16'd1230, 16'd18317, 16'd31151, 16'd33585, 16'd37284, 16'd12411, 16'd14657, 16'd13496}; // indx = 1411
    #10;
    addra = 32'd45184;
    dina = {96'd0, 16'd52645, 16'd47316, 16'd42972, 16'd29868, 16'd33241, 16'd876, 16'd6114, 16'd51700, 16'd14346, 16'd28225}; // indx = 1412
    #10;
    addra = 32'd45216;
    dina = {96'd0, 16'd55903, 16'd52501, 16'd26766, 16'd26437, 16'd4427, 16'd9229, 16'd44581, 16'd62981, 16'd25854, 16'd14693}; // indx = 1413
    #10;
    addra = 32'd45248;
    dina = {96'd0, 16'd59025, 16'd40318, 16'd36458, 16'd61894, 16'd23188, 16'd34136, 16'd32440, 16'd49257, 16'd19350, 16'd31936}; // indx = 1414
    #10;
    addra = 32'd45280;
    dina = {96'd0, 16'd33098, 16'd34603, 16'd32368, 16'd15980, 16'd28618, 16'd2659, 16'd13767, 16'd45669, 16'd33725, 16'd54175}; // indx = 1415
    #10;
    addra = 32'd45312;
    dina = {96'd0, 16'd35275, 16'd39653, 16'd32004, 16'd17322, 16'd55298, 16'd12241, 16'd47087, 16'd23288, 16'd15555, 16'd18525}; // indx = 1416
    #10;
    addra = 32'd45344;
    dina = {96'd0, 16'd24212, 16'd47599, 16'd39569, 16'd12321, 16'd13689, 16'd31033, 16'd31292, 16'd57817, 16'd40593, 16'd42150}; // indx = 1417
    #10;
    addra = 32'd45376;
    dina = {96'd0, 16'd52482, 16'd20146, 16'd44675, 16'd19541, 16'd65254, 16'd17606, 16'd39413, 16'd41122, 16'd35683, 16'd55408}; // indx = 1418
    #10;
    addra = 32'd45408;
    dina = {96'd0, 16'd7132, 16'd17551, 16'd17704, 16'd12997, 16'd25591, 16'd60680, 16'd57396, 16'd14628, 16'd25987, 16'd46485}; // indx = 1419
    #10;
    addra = 32'd45440;
    dina = {96'd0, 16'd32888, 16'd50612, 16'd29680, 16'd25873, 16'd28216, 16'd10654, 16'd47364, 16'd19130, 16'd4925, 16'd52941}; // indx = 1420
    #10;
    addra = 32'd45472;
    dina = {96'd0, 16'd49706, 16'd63249, 16'd14223, 16'd11467, 16'd60311, 16'd51904, 16'd15399, 16'd9738, 16'd24979, 16'd15845}; // indx = 1421
    #10;
    addra = 32'd45504;
    dina = {96'd0, 16'd24367, 16'd16801, 16'd19675, 16'd51358, 16'd3307, 16'd52721, 16'd24391, 16'd32411, 16'd7329, 16'd8762}; // indx = 1422
    #10;
    addra = 32'd45536;
    dina = {96'd0, 16'd43673, 16'd32519, 16'd33775, 16'd33220, 16'd23695, 16'd42171, 16'd55153, 16'd59120, 16'd26275, 16'd58506}; // indx = 1423
    #10;
    addra = 32'd45568;
    dina = {96'd0, 16'd25247, 16'd51657, 16'd64656, 16'd58879, 16'd46073, 16'd18875, 16'd21757, 16'd31543, 16'd49574, 16'd11940}; // indx = 1424
    #10;
    addra = 32'd45600;
    dina = {96'd0, 16'd47269, 16'd35249, 16'd48179, 16'd29993, 16'd34824, 16'd36952, 16'd51530, 16'd28226, 16'd48545, 16'd50485}; // indx = 1425
    #10;
    addra = 32'd45632;
    dina = {96'd0, 16'd8967, 16'd18702, 16'd24791, 16'd47821, 16'd58036, 16'd28807, 16'd16843, 16'd17144, 16'd48161, 16'd50490}; // indx = 1426
    #10;
    addra = 32'd45664;
    dina = {96'd0, 16'd16756, 16'd52361, 16'd55950, 16'd54164, 16'd26262, 16'd32582, 16'd44578, 16'd34926, 16'd13047, 16'd16209}; // indx = 1427
    #10;
    addra = 32'd45696;
    dina = {96'd0, 16'd54709, 16'd25007, 16'd22726, 16'd10321, 16'd43535, 16'd39029, 16'd36636, 16'd39031, 16'd62965, 16'd3982}; // indx = 1428
    #10;
    addra = 32'd45728;
    dina = {96'd0, 16'd52817, 16'd45427, 16'd54766, 16'd735, 16'd15451, 16'd8164, 16'd17716, 16'd8648, 16'd32643, 16'd45921}; // indx = 1429
    #10;
    addra = 32'd45760;
    dina = {96'd0, 16'd78, 16'd28723, 16'd58606, 16'd63224, 16'd58815, 16'd60724, 16'd27223, 16'd12168, 16'd51256, 16'd22059}; // indx = 1430
    #10;
    addra = 32'd45792;
    dina = {96'd0, 16'd32603, 16'd61585, 16'd31166, 16'd13687, 16'd55247, 16'd749, 16'd60997, 16'd34108, 16'd29282, 16'd30000}; // indx = 1431
    #10;
    addra = 32'd45824;
    dina = {96'd0, 16'd53163, 16'd62910, 16'd24041, 16'd32685, 16'd32897, 16'd50365, 16'd53545, 16'd44017, 16'd33146, 16'd5191}; // indx = 1432
    #10;
    addra = 32'd45856;
    dina = {96'd0, 16'd47529, 16'd38820, 16'd10131, 16'd57047, 16'd47792, 16'd41053, 16'd16391, 16'd57188, 16'd43911, 16'd29244}; // indx = 1433
    #10;
    addra = 32'd45888;
    dina = {96'd0, 16'd24468, 16'd58063, 16'd32410, 16'd46633, 16'd50103, 16'd26064, 16'd39303, 16'd13679, 16'd9064, 16'd53214}; // indx = 1434
    #10;
    addra = 32'd45920;
    dina = {96'd0, 16'd2935, 16'd60038, 16'd51429, 16'd37429, 16'd51292, 16'd20114, 16'd34132, 16'd1707, 16'd34596, 16'd20224}; // indx = 1435
    #10;
    addra = 32'd45952;
    dina = {96'd0, 16'd60762, 16'd34464, 16'd50583, 16'd50032, 16'd27017, 16'd63212, 16'd62996, 16'd38864, 16'd28761, 16'd30927}; // indx = 1436
    #10;
    addra = 32'd45984;
    dina = {96'd0, 16'd48050, 16'd57380, 16'd30544, 16'd29026, 16'd14567, 16'd25377, 16'd23728, 16'd39805, 16'd16617, 16'd44478}; // indx = 1437
    #10;
    addra = 32'd46016;
    dina = {96'd0, 16'd50418, 16'd42756, 16'd27443, 16'd17927, 16'd34481, 16'd53186, 16'd58025, 16'd5151, 16'd52270, 16'd30269}; // indx = 1438
    #10;
    addra = 32'd46048;
    dina = {96'd0, 16'd2192, 16'd33454, 16'd56678, 16'd8078, 16'd63005, 16'd61748, 16'd62367, 16'd31376, 16'd1460, 16'd53529}; // indx = 1439
    #10;
    addra = 32'd46080;
    dina = {96'd0, 16'd23294, 16'd64150, 16'd51946, 16'd62164, 16'd26960, 16'd48218, 16'd1735, 16'd20343, 16'd49637, 16'd35889}; // indx = 1440
    #10;
    addra = 32'd46112;
    dina = {96'd0, 16'd19067, 16'd21747, 16'd57216, 16'd1752, 16'd14856, 16'd30681, 16'd21758, 16'd44809, 16'd65504, 16'd52159}; // indx = 1441
    #10;
    addra = 32'd46144;
    dina = {96'd0, 16'd23033, 16'd60733, 16'd12038, 16'd11630, 16'd23424, 16'd37350, 16'd63057, 16'd62123, 16'd13980, 16'd16685}; // indx = 1442
    #10;
    addra = 32'd46176;
    dina = {96'd0, 16'd21870, 16'd38642, 16'd40111, 16'd14878, 16'd47047, 16'd33325, 16'd39385, 16'd46834, 16'd18042, 16'd25822}; // indx = 1443
    #10;
    addra = 32'd46208;
    dina = {96'd0, 16'd13122, 16'd44994, 16'd5007, 16'd41057, 16'd39423, 16'd63147, 16'd58356, 16'd55705, 16'd16985, 16'd6559}; // indx = 1444
    #10;
    addra = 32'd46240;
    dina = {96'd0, 16'd19868, 16'd40865, 16'd34067, 16'd12029, 16'd30783, 16'd39587, 16'd61036, 16'd45001, 16'd42661, 16'd19391}; // indx = 1445
    #10;
    addra = 32'd46272;
    dina = {96'd0, 16'd10785, 16'd33972, 16'd29712, 16'd33678, 16'd50607, 16'd17496, 16'd31945, 16'd30166, 16'd37953, 16'd3048}; // indx = 1446
    #10;
    addra = 32'd46304;
    dina = {96'd0, 16'd64546, 16'd41043, 16'd1994, 16'd25384, 16'd41917, 16'd57924, 16'd35319, 16'd13328, 16'd40855, 16'd55655}; // indx = 1447
    #10;
    addra = 32'd46336;
    dina = {96'd0, 16'd32732, 16'd6469, 16'd29549, 16'd26133, 16'd60899, 16'd18165, 16'd19501, 16'd44023, 16'd16298, 16'd24593}; // indx = 1448
    #10;
    addra = 32'd46368;
    dina = {96'd0, 16'd52621, 16'd27888, 16'd1059, 16'd27984, 16'd42066, 16'd49482, 16'd14206, 16'd51347, 16'd55003, 16'd58927}; // indx = 1449
    #10;
    addra = 32'd46400;
    dina = {96'd0, 16'd57762, 16'd59488, 16'd57250, 16'd37670, 16'd14448, 16'd39793, 16'd38007, 16'd48240, 16'd42945, 16'd25985}; // indx = 1450
    #10;
    addra = 32'd46432;
    dina = {96'd0, 16'd58138, 16'd264, 16'd24533, 16'd24858, 16'd42709, 16'd8003, 16'd33535, 16'd18868, 16'd44533, 16'd24786}; // indx = 1451
    #10;
    addra = 32'd46464;
    dina = {96'd0, 16'd6845, 16'd33908, 16'd45285, 16'd34950, 16'd11495, 16'd51861, 16'd60898, 16'd13865, 16'd20492, 16'd14836}; // indx = 1452
    #10;
    addra = 32'd46496;
    dina = {96'd0, 16'd32915, 16'd54162, 16'd34809, 16'd33678, 16'd33375, 16'd32604, 16'd19748, 16'd11756, 16'd8344, 16'd41886}; // indx = 1453
    #10;
    addra = 32'd46528;
    dina = {96'd0, 16'd17017, 16'd32381, 16'd33617, 16'd32819, 16'd61984, 16'd5444, 16'd23320, 16'd32257, 16'd47638, 16'd37781}; // indx = 1454
    #10;
    addra = 32'd46560;
    dina = {96'd0, 16'd20102, 16'd60078, 16'd50771, 16'd37570, 16'd33332, 16'd6163, 16'd31449, 16'd34784, 16'd5235, 16'd26361}; // indx = 1455
    #10;
    addra = 32'd46592;
    dina = {96'd0, 16'd58566, 16'd21001, 16'd49418, 16'd31361, 16'd56173, 16'd47280, 16'd17966, 16'd40000, 16'd23777, 16'd65498}; // indx = 1456
    #10;
    addra = 32'd46624;
    dina = {96'd0, 16'd34200, 16'd60725, 16'd16633, 16'd65048, 16'd6101, 16'd65024, 16'd18889, 16'd33545, 16'd39506, 16'd30163}; // indx = 1457
    #10;
    addra = 32'd46656;
    dina = {96'd0, 16'd36148, 16'd33658, 16'd8369, 16'd63613, 16'd57582, 16'd23568, 16'd54787, 16'd11816, 16'd22046, 16'd16274}; // indx = 1458
    #10;
    addra = 32'd46688;
    dina = {96'd0, 16'd53455, 16'd1686, 16'd56771, 16'd465, 16'd31469, 16'd40783, 16'd37107, 16'd65096, 16'd15353, 16'd46798}; // indx = 1459
    #10;
    addra = 32'd46720;
    dina = {96'd0, 16'd38489, 16'd38537, 16'd35827, 16'd16027, 16'd50700, 16'd26377, 16'd48351, 16'd41710, 16'd22368, 16'd2319}; // indx = 1460
    #10;
    addra = 32'd46752;
    dina = {96'd0, 16'd39093, 16'd55756, 16'd34724, 16'd54368, 16'd37354, 16'd11965, 16'd47069, 16'd5853, 16'd43900, 16'd5306}; // indx = 1461
    #10;
    addra = 32'd46784;
    dina = {96'd0, 16'd46968, 16'd57249, 16'd28075, 16'd9466, 16'd20385, 16'd56168, 16'd35979, 16'd54901, 16'd38246, 16'd31647}; // indx = 1462
    #10;
    addra = 32'd46816;
    dina = {96'd0, 16'd22615, 16'd63254, 16'd44627, 16'd23834, 16'd49318, 16'd13896, 16'd55409, 16'd27757, 16'd53701, 16'd7161}; // indx = 1463
    #10;
    addra = 32'd46848;
    dina = {96'd0, 16'd53587, 16'd37729, 16'd50717, 16'd38367, 16'd10086, 16'd61167, 16'd17681, 16'd63790, 16'd6214, 16'd51444}; // indx = 1464
    #10;
    addra = 32'd46880;
    dina = {96'd0, 16'd6735, 16'd39511, 16'd40080, 16'd26438, 16'd28279, 16'd41732, 16'd56180, 16'd17149, 16'd26866, 16'd60935}; // indx = 1465
    #10;
    addra = 32'd46912;
    dina = {96'd0, 16'd17610, 16'd44899, 16'd20973, 16'd9167, 16'd9483, 16'd19816, 16'd53895, 16'd49484, 16'd41601, 16'd31948}; // indx = 1466
    #10;
    addra = 32'd46944;
    dina = {96'd0, 16'd36004, 16'd38795, 16'd21843, 16'd27997, 16'd57575, 16'd25823, 16'd57258, 16'd5184, 16'd28989, 16'd12805}; // indx = 1467
    #10;
    addra = 32'd46976;
    dina = {96'd0, 16'd19422, 16'd51367, 16'd802, 16'd28878, 16'd793, 16'd23191, 16'd33474, 16'd53142, 16'd41533, 16'd40361}; // indx = 1468
    #10;
    addra = 32'd47008;
    dina = {96'd0, 16'd25714, 16'd53783, 16'd46664, 16'd18494, 16'd49849, 16'd17841, 16'd47717, 16'd4053, 16'd52493, 16'd36514}; // indx = 1469
    #10;
    addra = 32'd47040;
    dina = {96'd0, 16'd28978, 16'd43713, 16'd52565, 16'd30794, 16'd58218, 16'd55793, 16'd39632, 16'd58036, 16'd13680, 16'd9439}; // indx = 1470
    #10;
    addra = 32'd47072;
    dina = {96'd0, 16'd37486, 16'd48078, 16'd15353, 16'd61589, 16'd28914, 16'd36461, 16'd28906, 16'd25228, 16'd22642, 16'd20874}; // indx = 1471
    #10;
    addra = 32'd47104;
    dina = {96'd0, 16'd45453, 16'd52641, 16'd29563, 16'd64719, 16'd31878, 16'd36165, 16'd4559, 16'd24580, 16'd40027, 16'd58829}; // indx = 1472
    #10;
    addra = 32'd47136;
    dina = {96'd0, 16'd31797, 16'd11218, 16'd16812, 16'd21353, 16'd44176, 16'd54141, 16'd58887, 16'd49699, 16'd44074, 16'd3936}; // indx = 1473
    #10;
    addra = 32'd47168;
    dina = {96'd0, 16'd38313, 16'd8222, 16'd60551, 16'd41453, 16'd15324, 16'd29282, 16'd8045, 16'd38515, 16'd2678, 16'd3751}; // indx = 1474
    #10;
    addra = 32'd47200;
    dina = {96'd0, 16'd53358, 16'd57575, 16'd28356, 16'd2467, 16'd2784, 16'd31347, 16'd27503, 16'd5785, 16'd23115, 16'd58097}; // indx = 1475
    #10;
    addra = 32'd47232;
    dina = {96'd0, 16'd21818, 16'd21959, 16'd55436, 16'd40473, 16'd43894, 16'd43786, 16'd35661, 16'd51806, 16'd28425, 16'd18602}; // indx = 1476
    #10;
    addra = 32'd47264;
    dina = {96'd0, 16'd48780, 16'd26953, 16'd64609, 16'd24257, 16'd62689, 16'd53404, 16'd55201, 16'd22950, 16'd29196, 16'd46528}; // indx = 1477
    #10;
    addra = 32'd47296;
    dina = {96'd0, 16'd38389, 16'd38537, 16'd23122, 16'd56430, 16'd50618, 16'd58126, 16'd46213, 16'd27347, 16'd16117, 16'd55771}; // indx = 1478
    #10;
    addra = 32'd47328;
    dina = {96'd0, 16'd18105, 16'd566, 16'd53114, 16'd55867, 16'd54177, 16'd7570, 16'd58670, 16'd18997, 16'd50570, 16'd46955}; // indx = 1479
    #10;
    addra = 32'd47360;
    dina = {96'd0, 16'd21031, 16'd22575, 16'd59674, 16'd19765, 16'd62324, 16'd50975, 16'd65248, 16'd58323, 16'd28454, 16'd369}; // indx = 1480
    #10;
    addra = 32'd47392;
    dina = {96'd0, 16'd64493, 16'd986, 16'd59300, 16'd59137, 16'd52516, 16'd37103, 16'd1754, 16'd20358, 16'd64442, 16'd4338}; // indx = 1481
    #10;
    addra = 32'd47424;
    dina = {96'd0, 16'd57052, 16'd63530, 16'd47174, 16'd46064, 16'd46623, 16'd57362, 16'd38577, 16'd46697, 16'd1140, 16'd32135}; // indx = 1482
    #10;
    addra = 32'd47456;
    dina = {96'd0, 16'd57069, 16'd29403, 16'd8345, 16'd7953, 16'd23008, 16'd13924, 16'd19592, 16'd28210, 16'd11168, 16'd65073}; // indx = 1483
    #10;
    addra = 32'd47488;
    dina = {96'd0, 16'd29995, 16'd44691, 16'd19959, 16'd51249, 16'd58615, 16'd47298, 16'd21997, 16'd45475, 16'd19607, 16'd44938}; // indx = 1484
    #10;
    addra = 32'd47520;
    dina = {96'd0, 16'd15519, 16'd10544, 16'd36791, 16'd5983, 16'd57856, 16'd26257, 16'd1921, 16'd20639, 16'd58353, 16'd600}; // indx = 1485
    #10;
    addra = 32'd47552;
    dina = {96'd0, 16'd44989, 16'd32809, 16'd64763, 16'd34419, 16'd25834, 16'd107, 16'd59975, 16'd39878, 16'd14937, 16'd40601}; // indx = 1486
    #10;
    addra = 32'd47584;
    dina = {96'd0, 16'd65321, 16'd34532, 16'd10384, 16'd52667, 16'd9501, 16'd26914, 16'd13024, 16'd14047, 16'd30167, 16'd34262}; // indx = 1487
    #10;
    addra = 32'd47616;
    dina = {96'd0, 16'd25624, 16'd20130, 16'd19532, 16'd60716, 16'd1012, 16'd60732, 16'd63148, 16'd13066, 16'd34008, 16'd42413}; // indx = 1488
    #10;
    addra = 32'd47648;
    dina = {96'd0, 16'd42371, 16'd31537, 16'd37772, 16'd57543, 16'd53448, 16'd25686, 16'd30255, 16'd59409, 16'd24175, 16'd19954}; // indx = 1489
    #10;
    addra = 32'd47680;
    dina = {96'd0, 16'd4832, 16'd28952, 16'd29150, 16'd62181, 16'd8919, 16'd48399, 16'd17733, 16'd28116, 16'd59012, 16'd31374}; // indx = 1490
    #10;
    addra = 32'd47712;
    dina = {96'd0, 16'd41426, 16'd457, 16'd58242, 16'd29613, 16'd59180, 16'd25676, 16'd46492, 16'd21278, 16'd10530, 16'd61399}; // indx = 1491
    #10;
    addra = 32'd47744;
    dina = {96'd0, 16'd21086, 16'd23775, 16'd963, 16'd37325, 16'd51990, 16'd46218, 16'd10917, 16'd28637, 16'd22822, 16'd46206}; // indx = 1492
    #10;
    addra = 32'd47776;
    dina = {96'd0, 16'd3847, 16'd25015, 16'd1577, 16'd11675, 16'd14815, 16'd2880, 16'd22820, 16'd30253, 16'd8393, 16'd44920}; // indx = 1493
    #10;
    addra = 32'd47808;
    dina = {96'd0, 16'd37968, 16'd36498, 16'd60998, 16'd35274, 16'd45448, 16'd13546, 16'd60072, 16'd18153, 16'd34978, 16'd7836}; // indx = 1494
    #10;
    addra = 32'd47840;
    dina = {96'd0, 16'd48182, 16'd47060, 16'd48470, 16'd44886, 16'd50069, 16'd23713, 16'd665, 16'd844, 16'd20301, 16'd26235}; // indx = 1495
    #10;
    addra = 32'd47872;
    dina = {96'd0, 16'd43559, 16'd28824, 16'd7279, 16'd61336, 16'd31826, 16'd41262, 16'd20983, 16'd31987, 16'd21137, 16'd34954}; // indx = 1496
    #10;
    addra = 32'd47904;
    dina = {96'd0, 16'd26732, 16'd44796, 16'd39115, 16'd36412, 16'd23091, 16'd33247, 16'd24125, 16'd31564, 16'd33130, 16'd60517}; // indx = 1497
    #10;
    addra = 32'd47936;
    dina = {96'd0, 16'd20176, 16'd43173, 16'd47908, 16'd20002, 16'd62465, 16'd63190, 16'd39385, 16'd23015, 16'd303, 16'd4255}; // indx = 1498
    #10;
    addra = 32'd47968;
    dina = {96'd0, 16'd52895, 16'd9262, 16'd25304, 16'd1434, 16'd9863, 16'd19275, 16'd56007, 16'd42558, 16'd62771, 16'd9354}; // indx = 1499
    #10;
    addra = 32'd48000;
    dina = {96'd0, 16'd65011, 16'd12235, 16'd62522, 16'd24583, 16'd48197, 16'd55308, 16'd58588, 16'd28134, 16'd28162, 16'd46146}; // indx = 1500
    #10;
    addra = 32'd48032;
    dina = {96'd0, 16'd28034, 16'd64340, 16'd5006, 16'd30814, 16'd50435, 16'd42915, 16'd62466, 16'd46988, 16'd17457, 16'd37763}; // indx = 1501
    #10;
    addra = 32'd48064;
    dina = {96'd0, 16'd18187, 16'd16225, 16'd56645, 16'd30322, 16'd34198, 16'd40861, 16'd33200, 16'd15886, 16'd4856, 16'd62526}; // indx = 1502
    #10;
    addra = 32'd48096;
    dina = {96'd0, 16'd4831, 16'd16867, 16'd36518, 16'd52064, 16'd23643, 16'd41792, 16'd31900, 16'd25721, 16'd56127, 16'd63776}; // indx = 1503
    #10;
    addra = 32'd48128;
    dina = {96'd0, 16'd53399, 16'd34198, 16'd51980, 16'd10522, 16'd45639, 16'd19220, 16'd35526, 16'd34896, 16'd21235, 16'd55515}; // indx = 1504
    #10;
    addra = 32'd48160;
    dina = {96'd0, 16'd4561, 16'd21160, 16'd6832, 16'd14126, 16'd3549, 16'd42976, 16'd23866, 16'd56519, 16'd3847, 16'd34033}; // indx = 1505
    #10;
    addra = 32'd48192;
    dina = {96'd0, 16'd34095, 16'd10139, 16'd23041, 16'd50368, 16'd45518, 16'd10024, 16'd29027, 16'd24955, 16'd2506, 16'd18952}; // indx = 1506
    #10;
    addra = 32'd48224;
    dina = {96'd0, 16'd4140, 16'd31967, 16'd55361, 16'd6179, 16'd2417, 16'd19322, 16'd13983, 16'd53818, 16'd33226, 16'd53187}; // indx = 1507
    #10;
    addra = 32'd48256;
    dina = {96'd0, 16'd39655, 16'd25162, 16'd6528, 16'd2521, 16'd56394, 16'd37725, 16'd15452, 16'd1639, 16'd63240, 16'd29248}; // indx = 1508
    #10;
    addra = 32'd48288;
    dina = {96'd0, 16'd27362, 16'd13465, 16'd9336, 16'd51294, 16'd33394, 16'd59796, 16'd59149, 16'd63262, 16'd22537, 16'd21916}; // indx = 1509
    #10;
    addra = 32'd48320;
    dina = {96'd0, 16'd5419, 16'd38789, 16'd53653, 16'd20401, 16'd18220, 16'd56367, 16'd29377, 16'd46713, 16'd21212, 16'd2493}; // indx = 1510
    #10;
    addra = 32'd48352;
    dina = {96'd0, 16'd17368, 16'd29258, 16'd26634, 16'd21012, 16'd38078, 16'd22050, 16'd51839, 16'd22119, 16'd41852, 16'd45359}; // indx = 1511
    #10;
    addra = 32'd48384;
    dina = {96'd0, 16'd13953, 16'd51338, 16'd38860, 16'd58430, 16'd40191, 16'd22623, 16'd33733, 16'd6403, 16'd47111, 16'd7897}; // indx = 1512
    #10;
    addra = 32'd48416;
    dina = {96'd0, 16'd3326, 16'd12182, 16'd14385, 16'd8080, 16'd16983, 16'd11535, 16'd51498, 16'd2341, 16'd63630, 16'd43205}; // indx = 1513
    #10;
    addra = 32'd48448;
    dina = {96'd0, 16'd19916, 16'd4622, 16'd7721, 16'd10194, 16'd1577, 16'd5192, 16'd18933, 16'd5829, 16'd13405, 16'd64393}; // indx = 1514
    #10;
    addra = 32'd48480;
    dina = {96'd0, 16'd43396, 16'd32472, 16'd22333, 16'd45497, 16'd21580, 16'd54100, 16'd40958, 16'd3595, 16'd3630, 16'd34392}; // indx = 1515
    #10;
    addra = 32'd48512;
    dina = {96'd0, 16'd62783, 16'd31269, 16'd29459, 16'd24394, 16'd22630, 16'd47050, 16'd60497, 16'd22488, 16'd53239, 16'd27151}; // indx = 1516
    #10;
    addra = 32'd48544;
    dina = {96'd0, 16'd63938, 16'd40909, 16'd37340, 16'd32869, 16'd7215, 16'd49176, 16'd33049, 16'd19955, 16'd45294, 16'd25929}; // indx = 1517
    #10;
    addra = 32'd48576;
    dina = {96'd0, 16'd41962, 16'd5877, 16'd48532, 16'd49757, 16'd4633, 16'd418, 16'd2715, 16'd31566, 16'd19284, 16'd45723}; // indx = 1518
    #10;
    addra = 32'd48608;
    dina = {96'd0, 16'd56046, 16'd55638, 16'd33966, 16'd34688, 16'd8724, 16'd16839, 16'd28197, 16'd30010, 16'd42677, 16'd60340}; // indx = 1519
    #10;
    addra = 32'd48640;
    dina = {96'd0, 16'd43075, 16'd5639, 16'd51114, 16'd27949, 16'd11207, 16'd49753, 16'd22716, 16'd32936, 16'd27046, 16'd44754}; // indx = 1520
    #10;
    addra = 32'd48672;
    dina = {96'd0, 16'd60102, 16'd50677, 16'd63832, 16'd8841, 16'd47444, 16'd29073, 16'd45768, 16'd60342, 16'd30930, 16'd27272}; // indx = 1521
    #10;
    addra = 32'd48704;
    dina = {96'd0, 16'd50752, 16'd50549, 16'd6963, 16'd37139, 16'd61058, 16'd8852, 16'd21900, 16'd2272, 16'd63650, 16'd3562}; // indx = 1522
    #10;
    addra = 32'd48736;
    dina = {96'd0, 16'd23542, 16'd18689, 16'd63811, 16'd64820, 16'd30191, 16'd22373, 16'd61697, 16'd19579, 16'd7194, 16'd38308}; // indx = 1523
    #10;
    addra = 32'd48768;
    dina = {96'd0, 16'd20468, 16'd13084, 16'd38210, 16'd19591, 16'd7385, 16'd13952, 16'd17246, 16'd58429, 16'd59819, 16'd27691}; // indx = 1524
    #10;
    addra = 32'd48800;
    dina = {96'd0, 16'd11239, 16'd29940, 16'd25165, 16'd12575, 16'd43620, 16'd14971, 16'd145, 16'd22071, 16'd10360, 16'd64945}; // indx = 1525
    #10;
    addra = 32'd48832;
    dina = {96'd0, 16'd1829, 16'd20666, 16'd18625, 16'd1056, 16'd46788, 16'd61425, 16'd4286, 16'd56974, 16'd49823, 16'd43721}; // indx = 1526
    #10;
    addra = 32'd48864;
    dina = {96'd0, 16'd16183, 16'd16625, 16'd2493, 16'd4525, 16'd18520, 16'd36133, 16'd21783, 16'd55829, 16'd37405, 16'd20049}; // indx = 1527
    #10;
    addra = 32'd48896;
    dina = {96'd0, 16'd54250, 16'd34016, 16'd15416, 16'd31574, 16'd19794, 16'd7322, 16'd42414, 16'd30965, 16'd9591, 16'd48581}; // indx = 1528
    #10;
    addra = 32'd48928;
    dina = {96'd0, 16'd51210, 16'd57100, 16'd56260, 16'd28865, 16'd7134, 16'd3859, 16'd1627, 16'd499, 16'd6733, 16'd32215}; // indx = 1529
    #10;
    addra = 32'd48960;
    dina = {96'd0, 16'd926, 16'd46906, 16'd60007, 16'd18069, 16'd38989, 16'd7676, 16'd39902, 16'd12198, 16'd41513, 16'd12799}; // indx = 1530
    #10;
    addra = 32'd48992;
    dina = {96'd0, 16'd37476, 16'd13170, 16'd19770, 16'd52043, 16'd18475, 16'd1603, 16'd28942, 16'd65269, 16'd50919, 16'd45220}; // indx = 1531
    #10;
    addra = 32'd49024;
    dina = {96'd0, 16'd56679, 16'd12808, 16'd3604, 16'd43444, 16'd48334, 16'd41934, 16'd34495, 16'd38724, 16'd6140, 16'd65036}; // indx = 1532
    #10;
    addra = 32'd49056;
    dina = {96'd0, 16'd38576, 16'd58281, 16'd37401, 16'd52812, 16'd59107, 16'd4226, 16'd18017, 16'd32235, 16'd4265, 16'd23583}; // indx = 1533
    #10;
    addra = 32'd49088;
    dina = {96'd0, 16'd56152, 16'd61646, 16'd64783, 16'd56430, 16'd32572, 16'd59822, 16'd63165, 16'd22108, 16'd60558, 16'd5798}; // indx = 1534
    #10;
    addra = 32'd49120;
    dina = {96'd0, 16'd34251, 16'd55835, 16'd39037, 16'd12497, 16'd37886, 16'd57720, 16'd25886, 16'd48073, 16'd22538, 16'd52144}; // indx = 1535
    #10;
    addra = 32'd49152;
    dina = {96'd0, 16'd65356, 16'd60171, 16'd10417, 16'd37107, 16'd28424, 16'd60529, 16'd1026, 16'd35110, 16'd42956, 16'd47922}; // indx = 1536
    #10;
    addra = 32'd49184;
    dina = {96'd0, 16'd37349, 16'd19482, 16'd56585, 16'd45904, 16'd15677, 16'd26995, 16'd12158, 16'd58545, 16'd55994, 16'd12196}; // indx = 1537
    #10;
    addra = 32'd49216;
    dina = {96'd0, 16'd55691, 16'd18374, 16'd53916, 16'd9931, 16'd11918, 16'd61300, 16'd34085, 16'd52786, 16'd56940, 16'd41356}; // indx = 1538
    #10;
    addra = 32'd49248;
    dina = {96'd0, 16'd23985, 16'd30630, 16'd34205, 16'd21433, 16'd9637, 16'd10765, 16'd31993, 16'd23550, 16'd44054, 16'd37738}; // indx = 1539
    #10;
    addra = 32'd49280;
    dina = {96'd0, 16'd21794, 16'd13039, 16'd31285, 16'd57093, 16'd55905, 16'd35533, 16'd1604, 16'd9096, 16'd6947, 16'd19342}; // indx = 1540
    #10;
    addra = 32'd49312;
    dina = {96'd0, 16'd7100, 16'd47604, 16'd59132, 16'd5563, 16'd34451, 16'd33354, 16'd27859, 16'd42956, 16'd58360, 16'd43430}; // indx = 1541
    #10;
    addra = 32'd49344;
    dina = {96'd0, 16'd10420, 16'd54040, 16'd2352, 16'd4107, 16'd19309, 16'd39604, 16'd12920, 16'd60655, 16'd10672, 16'd34171}; // indx = 1542
    #10;
    addra = 32'd49376;
    dina = {96'd0, 16'd56240, 16'd27628, 16'd33376, 16'd43252, 16'd36854, 16'd2780, 16'd16048, 16'd9671, 16'd51594, 16'd47030}; // indx = 1543
    #10;
    addra = 32'd49408;
    dina = {96'd0, 16'd53126, 16'd5626, 16'd50000, 16'd40788, 16'd8940, 16'd3340, 16'd64564, 16'd39844, 16'd20039, 16'd946}; // indx = 1544
    #10;
    addra = 32'd49440;
    dina = {96'd0, 16'd11809, 16'd5856, 16'd60886, 16'd43054, 16'd58489, 16'd37583, 16'd2504, 16'd52692, 16'd58445, 16'd8742}; // indx = 1545
    #10;
    addra = 32'd49472;
    dina = {96'd0, 16'd52205, 16'd23134, 16'd30987, 16'd45671, 16'd17585, 16'd22451, 16'd8969, 16'd52350, 16'd25136, 16'd58866}; // indx = 1546
    #10;
    addra = 32'd49504;
    dina = {96'd0, 16'd25735, 16'd53510, 16'd52399, 16'd10093, 16'd45275, 16'd53771, 16'd34463, 16'd37623, 16'd167, 16'd62311}; // indx = 1547
    #10;
    addra = 32'd49536;
    dina = {96'd0, 16'd18508, 16'd19882, 16'd63088, 16'd36587, 16'd27739, 16'd60381, 16'd57489, 16'd17563, 16'd60225, 16'd5867}; // indx = 1548
    #10;
    addra = 32'd49568;
    dina = {96'd0, 16'd56548, 16'd12660, 16'd22070, 16'd43262, 16'd33563, 16'd42926, 16'd28702, 16'd43768, 16'd37364, 16'd21931}; // indx = 1549
    #10;
    addra = 32'd49600;
    dina = {96'd0, 16'd42818, 16'd51344, 16'd11416, 16'd58628, 16'd43579, 16'd65529, 16'd40996, 16'd2069, 16'd6698, 16'd53868}; // indx = 1550
    #10;
    addra = 32'd49632;
    dina = {96'd0, 16'd39692, 16'd59836, 16'd54616, 16'd64563, 16'd20584, 16'd17812, 16'd37443, 16'd46181, 16'd11346, 16'd3832}; // indx = 1551
    #10;
    addra = 32'd49664;
    dina = {96'd0, 16'd51718, 16'd34810, 16'd36354, 16'd17811, 16'd28876, 16'd21680, 16'd13681, 16'd56408, 16'd27177, 16'd6369}; // indx = 1552
    #10;
    addra = 32'd49696;
    dina = {96'd0, 16'd29141, 16'd52070, 16'd34467, 16'd37444, 16'd39313, 16'd725, 16'd27911, 16'd36389, 16'd30937, 16'd64784}; // indx = 1553
    #10;
    addra = 32'd49728;
    dina = {96'd0, 16'd45363, 16'd55652, 16'd59379, 16'd44963, 16'd47347, 16'd60555, 16'd40171, 16'd63273, 16'd53040, 16'd62751}; // indx = 1554
    #10;
    addra = 32'd49760;
    dina = {96'd0, 16'd58188, 16'd2819, 16'd60242, 16'd64117, 16'd9246, 16'd58014, 16'd43669, 16'd45664, 16'd17360, 16'd34777}; // indx = 1555
    #10;
    addra = 32'd49792;
    dina = {96'd0, 16'd28823, 16'd44713, 16'd40889, 16'd49407, 16'd31233, 16'd16307, 16'd6905, 16'd49153, 16'd46613, 16'd60973}; // indx = 1556
    #10;
    addra = 32'd49824;
    dina = {96'd0, 16'd36051, 16'd4384, 16'd55385, 16'd50241, 16'd52493, 16'd35524, 16'd16727, 16'd16906, 16'd37457, 16'd58640}; // indx = 1557
    #10;
    addra = 32'd49856;
    dina = {96'd0, 16'd32029, 16'd10488, 16'd60408, 16'd35780, 16'd20215, 16'd46448, 16'd54128, 16'd37276, 16'd54259, 16'd24734}; // indx = 1558
    #10;
    addra = 32'd49888;
    dina = {96'd0, 16'd12338, 16'd12487, 16'd35859, 16'd64194, 16'd42022, 16'd57543, 16'd27729, 16'd7361, 16'd37405, 16'd28444}; // indx = 1559
    #10;
    addra = 32'd49920;
    dina = {96'd0, 16'd9450, 16'd31166, 16'd32610, 16'd43101, 16'd62847, 16'd46774, 16'd17938, 16'd33083, 16'd53056, 16'd41049}; // indx = 1560
    #10;
    addra = 32'd49952;
    dina = {96'd0, 16'd35207, 16'd32304, 16'd44275, 16'd19476, 16'd8123, 16'd5205, 16'd22539, 16'd59929, 16'd45446, 16'd62179}; // indx = 1561
    #10;
    addra = 32'd49984;
    dina = {96'd0, 16'd35164, 16'd22, 16'd41421, 16'd24878, 16'd55457, 16'd45343, 16'd52778, 16'd42166, 16'd11950, 16'd6553}; // indx = 1562
    #10;
    addra = 32'd50016;
    dina = {96'd0, 16'd47701, 16'd12201, 16'd41149, 16'd31184, 16'd60287, 16'd7177, 16'd50983, 16'd44877, 16'd26865, 16'd49826}; // indx = 1563
    #10;
    addra = 32'd50048;
    dina = {96'd0, 16'd51098, 16'd34042, 16'd61956, 16'd10411, 16'd26172, 16'd52262, 16'd38541, 16'd24511, 16'd55826, 16'd17692}; // indx = 1564
    #10;
    addra = 32'd50080;
    dina = {96'd0, 16'd37333, 16'd28625, 16'd54860, 16'd10319, 16'd37759, 16'd14106, 16'd56666, 16'd29555, 16'd51300, 16'd57051}; // indx = 1565
    #10;
    addra = 32'd50112;
    dina = {96'd0, 16'd7734, 16'd32947, 16'd31394, 16'd1572, 16'd45969, 16'd59085, 16'd1476, 16'd20236, 16'd24905, 16'd63258}; // indx = 1566
    #10;
    addra = 32'd50144;
    dina = {96'd0, 16'd32858, 16'd24415, 16'd47815, 16'd388, 16'd43127, 16'd63924, 16'd11835, 16'd18570, 16'd15746, 16'd39587}; // indx = 1567
    #10;
    addra = 32'd50176;
    dina = {96'd0, 16'd12437, 16'd59603, 16'd14178, 16'd6766, 16'd58457, 16'd27833, 16'd15175, 16'd24383, 16'd51801, 16'd35144}; // indx = 1568
    #10;
    addra = 32'd50208;
    dina = {96'd0, 16'd5423, 16'd44831, 16'd25866, 16'd19522, 16'd56199, 16'd14115, 16'd50163, 16'd29207, 16'd3512, 16'd33129}; // indx = 1569
    #10;
    addra = 32'd50240;
    dina = {96'd0, 16'd1699, 16'd46467, 16'd37919, 16'd6107, 16'd3055, 16'd66, 16'd5430, 16'd26609, 16'd16472, 16'd59877}; // indx = 1570
    #10;
    addra = 32'd50272;
    dina = {96'd0, 16'd52094, 16'd38050, 16'd20091, 16'd57568, 16'd34121, 16'd34159, 16'd10685, 16'd15092, 16'd18601, 16'd49637}; // indx = 1571
    #10;
    addra = 32'd50304;
    dina = {96'd0, 16'd8655, 16'd5177, 16'd15382, 16'd36808, 16'd30435, 16'd27643, 16'd51740, 16'd34350, 16'd6480, 16'd17909}; // indx = 1572
    #10;
    addra = 32'd50336;
    dina = {96'd0, 16'd37671, 16'd57087, 16'd41172, 16'd32155, 16'd51183, 16'd50741, 16'd52835, 16'd35584, 16'd60632, 16'd44325}; // indx = 1573
    #10;
    addra = 32'd50368;
    dina = {96'd0, 16'd16104, 16'd25764, 16'd57535, 16'd30744, 16'd11204, 16'd41115, 16'd58071, 16'd59072, 16'd47156, 16'd13194}; // indx = 1574
    #10;
    addra = 32'd50400;
    dina = {96'd0, 16'd17366, 16'd9032, 16'd51134, 16'd23078, 16'd52078, 16'd12979, 16'd62430, 16'd38131, 16'd49235, 16'd4992}; // indx = 1575
    #10;
    addra = 32'd50432;
    dina = {96'd0, 16'd22477, 16'd52912, 16'd47937, 16'd54988, 16'd55067, 16'd31132, 16'd27490, 16'd34966, 16'd2927, 16'd13777}; // indx = 1576
    #10;
    addra = 32'd50464;
    dina = {96'd0, 16'd59680, 16'd55591, 16'd22757, 16'd7762, 16'd2479, 16'd4379, 16'd22358, 16'd45913, 16'd5641, 16'd23802}; // indx = 1577
    #10;
    addra = 32'd50496;
    dina = {96'd0, 16'd39782, 16'd50139, 16'd33552, 16'd57470, 16'd58344, 16'd12201, 16'd19168, 16'd40429, 16'd49367, 16'd27478}; // indx = 1578
    #10;
    addra = 32'd50528;
    dina = {96'd0, 16'd49572, 16'd24333, 16'd31354, 16'd4411, 16'd40959, 16'd25829, 16'd19515, 16'd65494, 16'd2886, 16'd777}; // indx = 1579
    #10;
    addra = 32'd50560;
    dina = {96'd0, 16'd64269, 16'd47614, 16'd8126, 16'd9632, 16'd44313, 16'd61462, 16'd7663, 16'd60682, 16'd10894, 16'd31305}; // indx = 1580
    #10;
    addra = 32'd50592;
    dina = {96'd0, 16'd31827, 16'd29136, 16'd62247, 16'd32889, 16'd60759, 16'd9723, 16'd58866, 16'd13423, 16'd63403, 16'd65201}; // indx = 1581
    #10;
    addra = 32'd50624;
    dina = {96'd0, 16'd53141, 16'd53649, 16'd21482, 16'd47794, 16'd25611, 16'd40400, 16'd46316, 16'd12519, 16'd31229, 16'd24029}; // indx = 1582
    #10;
    addra = 32'd50656;
    dina = {96'd0, 16'd55871, 16'd1856, 16'd18639, 16'd47720, 16'd64736, 16'd5269, 16'd31525, 16'd23863, 16'd41230, 16'd62641}; // indx = 1583
    #10;
    addra = 32'd50688;
    dina = {96'd0, 16'd10698, 16'd49020, 16'd13697, 16'd40136, 16'd60462, 16'd8951, 16'd4591, 16'd921, 16'd32840, 16'd65020}; // indx = 1584
    #10;
    addra = 32'd50720;
    dina = {96'd0, 16'd30048, 16'd24111, 16'd9434, 16'd62376, 16'd14680, 16'd29448, 16'd61452, 16'd25772, 16'd33132, 16'd15991}; // indx = 1585
    #10;
    addra = 32'd50752;
    dina = {96'd0, 16'd54744, 16'd26994, 16'd2182, 16'd57610, 16'd37859, 16'd24243, 16'd3291, 16'd64524, 16'd57458, 16'd63869}; // indx = 1586
    #10;
    addra = 32'd50784;
    dina = {96'd0, 16'd56096, 16'd14470, 16'd2652, 16'd37872, 16'd23766, 16'd14593, 16'd7174, 16'd15496, 16'd59804, 16'd41811}; // indx = 1587
    #10;
    addra = 32'd50816;
    dina = {96'd0, 16'd59612, 16'd28297, 16'd58742, 16'd51671, 16'd5399, 16'd64973, 16'd47066, 16'd49947, 16'd14352, 16'd43307}; // indx = 1588
    #10;
    addra = 32'd50848;
    dina = {96'd0, 16'd52445, 16'd3029, 16'd11673, 16'd34910, 16'd41437, 16'd24320, 16'd27779, 16'd44325, 16'd23607, 16'd61067}; // indx = 1589
    #10;
    addra = 32'd50880;
    dina = {96'd0, 16'd28510, 16'd9068, 16'd28280, 16'd1365, 16'd45612, 16'd40814, 16'd45172, 16'd10721, 16'd59706, 16'd34192}; // indx = 1590
    #10;
    addra = 32'd50912;
    dina = {96'd0, 16'd14285, 16'd26574, 16'd58838, 16'd35251, 16'd41289, 16'd5557, 16'd17235, 16'd29977, 16'd35454, 16'd22110}; // indx = 1591
    #10;
    addra = 32'd50944;
    dina = {96'd0, 16'd22451, 16'd33830, 16'd49711, 16'd18334, 16'd61510, 16'd20305, 16'd8459, 16'd44923, 16'd48209, 16'd35999}; // indx = 1592
    #10;
    addra = 32'd50976;
    dina = {96'd0, 16'd37091, 16'd27108, 16'd6754, 16'd64475, 16'd56235, 16'd24571, 16'd54250, 16'd3867, 16'd8449, 16'd24950}; // indx = 1593
    #10;
    addra = 32'd51008;
    dina = {96'd0, 16'd7225, 16'd885, 16'd17205, 16'd62183, 16'd39588, 16'd19736, 16'd35477, 16'd50101, 16'd9283, 16'd50367}; // indx = 1594
    #10;
    addra = 32'd51040;
    dina = {96'd0, 16'd1840, 16'd41410, 16'd33265, 16'd37502, 16'd21687, 16'd2829, 16'd34373, 16'd40032, 16'd7330, 16'd51065}; // indx = 1595
    #10;
    addra = 32'd51072;
    dina = {96'd0, 16'd53309, 16'd8266, 16'd52317, 16'd20367, 16'd12824, 16'd61008, 16'd11110, 16'd31618, 16'd30194, 16'd33548}; // indx = 1596
    #10;
    addra = 32'd51104;
    dina = {96'd0, 16'd15755, 16'd40082, 16'd12314, 16'd35723, 16'd61831, 16'd971, 16'd55459, 16'd4658, 16'd47995, 16'd6186}; // indx = 1597
    #10;
    addra = 32'd51136;
    dina = {96'd0, 16'd28515, 16'd40353, 16'd52661, 16'd57157, 16'd61913, 16'd23457, 16'd39563, 16'd43799, 16'd2977, 16'd44376}; // indx = 1598
    #10;
    addra = 32'd51168;
    dina = {96'd0, 16'd20984, 16'd60279, 16'd58155, 16'd9315, 16'd36490, 16'd44474, 16'd43079, 16'd51195, 16'd16160, 16'd43843}; // indx = 1599
    #10;
    addra = 32'd51200;
    dina = {96'd0, 16'd60519, 16'd46193, 16'd62284, 16'd9179, 16'd17790, 16'd36648, 16'd46650, 16'd3138, 16'd45606, 16'd8396}; // indx = 1600
    #10;
    addra = 32'd51232;
    dina = {96'd0, 16'd51439, 16'd36225, 16'd39439, 16'd56221, 16'd41580, 16'd59776, 16'd24310, 16'd5592, 16'd54315, 16'd8329}; // indx = 1601
    #10;
    addra = 32'd51264;
    dina = {96'd0, 16'd23575, 16'd59932, 16'd54610, 16'd42092, 16'd27167, 16'd28689, 16'd8805, 16'd12328, 16'd43232, 16'd335}; // indx = 1602
    #10;
    addra = 32'd51296;
    dina = {96'd0, 16'd45333, 16'd61025, 16'd35119, 16'd55550, 16'd50393, 16'd9194, 16'd55725, 16'd33224, 16'd697, 16'd60486}; // indx = 1603
    #10;
    addra = 32'd51328;
    dina = {96'd0, 16'd22791, 16'd13451, 16'd61265, 16'd24043, 16'd45090, 16'd37246, 16'd51233, 16'd46751, 16'd26278, 16'd36227}; // indx = 1604
    #10;
    addra = 32'd51360;
    dina = {96'd0, 16'd32374, 16'd31398, 16'd19494, 16'd39935, 16'd44618, 16'd43697, 16'd32179, 16'd37911, 16'd29650, 16'd51884}; // indx = 1605
    #10;
    addra = 32'd51392;
    dina = {96'd0, 16'd491, 16'd43901, 16'd10285, 16'd59200, 16'd37241, 16'd34927, 16'd26668, 16'd12329, 16'd27287, 16'd43977}; // indx = 1606
    #10;
    addra = 32'd51424;
    dina = {96'd0, 16'd29107, 16'd47324, 16'd2343, 16'd26259, 16'd521, 16'd8990, 16'd12084, 16'd54017, 16'd41401, 16'd31469}; // indx = 1607
    #10;
    addra = 32'd51456;
    dina = {96'd0, 16'd10046, 16'd4016, 16'd33020, 16'd24425, 16'd35584, 16'd22397, 16'd43976, 16'd46463, 16'd15597, 16'd43398}; // indx = 1608
    #10;
    addra = 32'd51488;
    dina = {96'd0, 16'd25413, 16'd13574, 16'd45637, 16'd12733, 16'd7085, 16'd54040, 16'd45649, 16'd26187, 16'd6372, 16'd53833}; // indx = 1609
    #10;
    addra = 32'd51520;
    dina = {96'd0, 16'd52521, 16'd38599, 16'd7527, 16'd9792, 16'd63622, 16'd8582, 16'd44027, 16'd34593, 16'd11856, 16'd51712}; // indx = 1610
    #10;
    addra = 32'd51552;
    dina = {96'd0, 16'd5020, 16'd16273, 16'd49054, 16'd58981, 16'd65121, 16'd4581, 16'd50037, 16'd20731, 16'd232, 16'd34563}; // indx = 1611
    #10;
    addra = 32'd51584;
    dina = {96'd0, 16'd56485, 16'd49365, 16'd15601, 16'd4042, 16'd28843, 16'd41758, 16'd58488, 16'd47750, 16'd40987, 16'd38289}; // indx = 1612
    #10;
    addra = 32'd51616;
    dina = {96'd0, 16'd33086, 16'd59995, 16'd46782, 16'd54702, 16'd33181, 16'd58271, 16'd52461, 16'd9238, 16'd11705, 16'd63874}; // indx = 1613
    #10;
    addra = 32'd51648;
    dina = {96'd0, 16'd8298, 16'd44711, 16'd47715, 16'd64679, 16'd51515, 16'd64433, 16'd3274, 16'd10191, 16'd31260, 16'd48080}; // indx = 1614
    #10;
    addra = 32'd51680;
    dina = {96'd0, 16'd57558, 16'd24178, 16'd10782, 16'd40883, 16'd52856, 16'd55130, 16'd13364, 16'd17000, 16'd49876, 16'd14095}; // indx = 1615
    #10;
    addra = 32'd51712;
    dina = {96'd0, 16'd46890, 16'd60352, 16'd11547, 16'd26586, 16'd16043, 16'd11686, 16'd1690, 16'd48913, 16'd54538, 16'd45699}; // indx = 1616
    #10;
    addra = 32'd51744;
    dina = {96'd0, 16'd37670, 16'd4022, 16'd51542, 16'd27615, 16'd9224, 16'd6467, 16'd11443, 16'd30943, 16'd15677, 16'd15458}; // indx = 1617
    #10;
    addra = 32'd51776;
    dina = {96'd0, 16'd18877, 16'd54510, 16'd43649, 16'd41864, 16'd39218, 16'd32838, 16'd45293, 16'd57405, 16'd2642, 16'd40404}; // indx = 1618
    #10;
    addra = 32'd51808;
    dina = {96'd0, 16'd5510, 16'd31751, 16'd27578, 16'd37036, 16'd28801, 16'd16818, 16'd59221, 16'd13831, 16'd42310, 16'd59931}; // indx = 1619
    #10;
    addra = 32'd51840;
    dina = {96'd0, 16'd18657, 16'd41010, 16'd59256, 16'd18216, 16'd21548, 16'd7367, 16'd6960, 16'd47045, 16'd58906, 16'd48711}; // indx = 1620
    #10;
    addra = 32'd51872;
    dina = {96'd0, 16'd39889, 16'd35059, 16'd2839, 16'd61437, 16'd18133, 16'd56149, 16'd34479, 16'd10048, 16'd33195, 16'd27859}; // indx = 1621
    #10;
    addra = 32'd51904;
    dina = {96'd0, 16'd9972, 16'd35254, 16'd11856, 16'd19631, 16'd18483, 16'd59474, 16'd30644, 16'd51688, 16'd62729, 16'd57750}; // indx = 1622
    #10;
    addra = 32'd51936;
    dina = {96'd0, 16'd40002, 16'd64497, 16'd31646, 16'd13970, 16'd43240, 16'd20638, 16'd22183, 16'd38919, 16'd1744, 16'd19178}; // indx = 1623
    #10;
    addra = 32'd51968;
    dina = {96'd0, 16'd7024, 16'd45782, 16'd41073, 16'd2171, 16'd57035, 16'd45780, 16'd10126, 16'd48040, 16'd36992, 16'd2929}; // indx = 1624
    #10;
    addra = 32'd52000;
    dina = {96'd0, 16'd31322, 16'd3541, 16'd27260, 16'd3022, 16'd4358, 16'd50731, 16'd30272, 16'd8779, 16'd65437, 16'd44200}; // indx = 1625
    #10;
    addra = 32'd52032;
    dina = {96'd0, 16'd48206, 16'd18824, 16'd46677, 16'd55550, 16'd47217, 16'd7536, 16'd5996, 16'd2535, 16'd37797, 16'd29676}; // indx = 1626
    #10;
    addra = 32'd52064;
    dina = {96'd0, 16'd55013, 16'd21167, 16'd31780, 16'd38049, 16'd39510, 16'd42459, 16'd50761, 16'd5042, 16'd19434, 16'd28021}; // indx = 1627
    #10;
    addra = 32'd52096;
    dina = {96'd0, 16'd25317, 16'd5302, 16'd61279, 16'd33698, 16'd32712, 16'd46916, 16'd21026, 16'd64972, 16'd3875, 16'd28874}; // indx = 1628
    #10;
    addra = 32'd52128;
    dina = {96'd0, 16'd18166, 16'd331, 16'd46804, 16'd35924, 16'd25094, 16'd17623, 16'd29786, 16'd20292, 16'd37484, 16'd29413}; // indx = 1629
    #10;
    addra = 32'd52160;
    dina = {96'd0, 16'd54377, 16'd15002, 16'd30956, 16'd58418, 16'd27756, 16'd18848, 16'd31018, 16'd58297, 16'd51138, 16'd53476}; // indx = 1630
    #10;
    addra = 32'd52192;
    dina = {96'd0, 16'd57147, 16'd18447, 16'd30861, 16'd1099, 16'd46001, 16'd37900, 16'd63630, 16'd39357, 16'd38251, 16'd12442}; // indx = 1631
    #10;
    addra = 32'd52224;
    dina = {96'd0, 16'd6239, 16'd52627, 16'd63664, 16'd9976, 16'd35181, 16'd15792, 16'd30972, 16'd52399, 16'd49427, 16'd34908}; // indx = 1632
    #10;
    addra = 32'd52256;
    dina = {96'd0, 16'd23477, 16'd52248, 16'd1282, 16'd47690, 16'd6032, 16'd18195, 16'd25182, 16'd39592, 16'd54476, 16'd34226}; // indx = 1633
    #10;
    addra = 32'd52288;
    dina = {96'd0, 16'd50930, 16'd52198, 16'd450, 16'd53426, 16'd51935, 16'd42581, 16'd51339, 16'd15469, 16'd36482, 16'd53306}; // indx = 1634
    #10;
    addra = 32'd52320;
    dina = {96'd0, 16'd31027, 16'd47670, 16'd61444, 16'd33909, 16'd59252, 16'd14306, 16'd5445, 16'd1141, 16'd60533, 16'd46467}; // indx = 1635
    #10;
    addra = 32'd52352;
    dina = {96'd0, 16'd56296, 16'd38468, 16'd5325, 16'd54061, 16'd29162, 16'd2831, 16'd9556, 16'd53867, 16'd19682, 16'd34853}; // indx = 1636
    #10;
    addra = 32'd52384;
    dina = {96'd0, 16'd41789, 16'd62368, 16'd57126, 16'd51185, 16'd31574, 16'd26580, 16'd56160, 16'd38063, 16'd16850, 16'd41401}; // indx = 1637
    #10;
    addra = 32'd52416;
    dina = {96'd0, 16'd22875, 16'd59340, 16'd48573, 16'd3338, 16'd25942, 16'd49948, 16'd47128, 16'd55487, 16'd29190, 16'd436}; // indx = 1638
    #10;
    addra = 32'd52448;
    dina = {96'd0, 16'd10575, 16'd45960, 16'd60695, 16'd36247, 16'd32605, 16'd60274, 16'd49746, 16'd6607, 16'd38620, 16'd38620}; // indx = 1639
    #10;
    addra = 32'd52480;
    dina = {96'd0, 16'd34375, 16'd47379, 16'd32005, 16'd41409, 16'd51593, 16'd3901, 16'd51474, 16'd45228, 16'd57056, 16'd33812}; // indx = 1640
    #10;
    addra = 32'd52512;
    dina = {96'd0, 16'd33989, 16'd9143, 16'd52381, 16'd50253, 16'd3732, 16'd8551, 16'd62005, 16'd40498, 16'd52099, 16'd22902}; // indx = 1641
    #10;
    addra = 32'd52544;
    dina = {96'd0, 16'd50050, 16'd56291, 16'd25141, 16'd20995, 16'd52869, 16'd6313, 16'd19399, 16'd60551, 16'd54877, 16'd44533}; // indx = 1642
    #10;
    addra = 32'd52576;
    dina = {96'd0, 16'd55831, 16'd7867, 16'd36345, 16'd9811, 16'd13561, 16'd55417, 16'd28350, 16'd61596, 16'd15997, 16'd21354}; // indx = 1643
    #10;
    addra = 32'd52608;
    dina = {96'd0, 16'd30845, 16'd31930, 16'd50927, 16'd36914, 16'd45305, 16'd63966, 16'd49346, 16'd26245, 16'd35690, 16'd18016}; // indx = 1644
    #10;
    addra = 32'd52640;
    dina = {96'd0, 16'd36423, 16'd25163, 16'd28090, 16'd9866, 16'd3121, 16'd19750, 16'd5712, 16'd50189, 16'd49796, 16'd1864}; // indx = 1645
    #10;
    addra = 32'd52672;
    dina = {96'd0, 16'd7553, 16'd27728, 16'd34791, 16'd43007, 16'd53289, 16'd54819, 16'd14902, 16'd60547, 16'd62203, 16'd17691}; // indx = 1646
    #10;
    addra = 32'd52704;
    dina = {96'd0, 16'd51786, 16'd21119, 16'd49790, 16'd55888, 16'd20648, 16'd7680, 16'd4527, 16'd27502, 16'd21034, 16'd11073}; // indx = 1647
    #10;
    addra = 32'd52736;
    dina = {96'd0, 16'd48860, 16'd45686, 16'd45472, 16'd25284, 16'd36922, 16'd29060, 16'd44081, 16'd40729, 16'd6900, 16'd28082}; // indx = 1648
    #10;
    addra = 32'd52768;
    dina = {96'd0, 16'd16730, 16'd17142, 16'd15598, 16'd62289, 16'd6235, 16'd25403, 16'd57221, 16'd21268, 16'd34340, 16'd22934}; // indx = 1649
    #10;
    addra = 32'd52800;
    dina = {96'd0, 16'd21527, 16'd9708, 16'd60504, 16'd46718, 16'd15923, 16'd26983, 16'd32998, 16'd46145, 16'd1710, 16'd12865}; // indx = 1650
    #10;
    addra = 32'd52832;
    dina = {96'd0, 16'd24931, 16'd63356, 16'd51526, 16'd53880, 16'd16593, 16'd35394, 16'd13728, 16'd15914, 16'd35934, 16'd3215}; // indx = 1651
    #10;
    addra = 32'd52864;
    dina = {96'd0, 16'd59060, 16'd65360, 16'd12237, 16'd5774, 16'd39011, 16'd8972, 16'd10269, 16'd42977, 16'd22156, 16'd33919}; // indx = 1652
    #10;
    addra = 32'd52896;
    dina = {96'd0, 16'd601, 16'd14698, 16'd48959, 16'd61042, 16'd52189, 16'd25556, 16'd58061, 16'd50740, 16'd63148, 16'd22923}; // indx = 1653
    #10;
    addra = 32'd52928;
    dina = {96'd0, 16'd40027, 16'd22189, 16'd54899, 16'd25395, 16'd11294, 16'd19762, 16'd37003, 16'd23719, 16'd22967, 16'd58693}; // indx = 1654
    #10;
    addra = 32'd52960;
    dina = {96'd0, 16'd44692, 16'd16794, 16'd61673, 16'd63769, 16'd16140, 16'd15537, 16'd30435, 16'd42215, 16'd23816, 16'd22659}; // indx = 1655
    #10;
    addra = 32'd52992;
    dina = {96'd0, 16'd35288, 16'd2270, 16'd9824, 16'd39002, 16'd2235, 16'd30949, 16'd26685, 16'd61134, 16'd52989, 16'd28628}; // indx = 1656
    #10;
    addra = 32'd53024;
    dina = {96'd0, 16'd58235, 16'd9699, 16'd59303, 16'd17566, 16'd29863, 16'd43996, 16'd13608, 16'd55566, 16'd34479, 16'd37364}; // indx = 1657
    #10;
    addra = 32'd53056;
    dina = {96'd0, 16'd50587, 16'd56616, 16'd35128, 16'd37204, 16'd34910, 16'd6491, 16'd33586, 16'd2533, 16'd56681, 16'd784}; // indx = 1658
    #10;
    addra = 32'd53088;
    dina = {96'd0, 16'd16826, 16'd14948, 16'd65221, 16'd33145, 16'd18160, 16'd24906, 16'd6204, 16'd30872, 16'd17401, 16'd18686}; // indx = 1659
    #10;
    addra = 32'd53120;
    dina = {96'd0, 16'd16991, 16'd2514, 16'd20158, 16'd52070, 16'd39847, 16'd56070, 16'd52960, 16'd60698, 16'd29122, 16'd61596}; // indx = 1660
    #10;
    addra = 32'd53152;
    dina = {96'd0, 16'd2291, 16'd33292, 16'd20576, 16'd31190, 16'd20502, 16'd28478, 16'd64183, 16'd19680, 16'd20689, 16'd42046}; // indx = 1661
    #10;
    addra = 32'd53184;
    dina = {96'd0, 16'd39249, 16'd18095, 16'd34022, 16'd245, 16'd7080, 16'd11284, 16'd6515, 16'd8845, 16'd19891, 16'd50337}; // indx = 1662
    #10;
    addra = 32'd53216;
    dina = {96'd0, 16'd38601, 16'd55895, 16'd40472, 16'd38786, 16'd41949, 16'd41866, 16'd47568, 16'd26670, 16'd62569, 16'd18115}; // indx = 1663
    #10;
    addra = 32'd53248;
    dina = {96'd0, 16'd26384, 16'd25519, 16'd60366, 16'd46783, 16'd44999, 16'd13138, 16'd42728, 16'd3317, 16'd9185, 16'd32378}; // indx = 1664
    #10;
    addra = 32'd53280;
    dina = {96'd0, 16'd8089, 16'd31767, 16'd46785, 16'd64999, 16'd18075, 16'd54024, 16'd26816, 16'd18972, 16'd43222, 16'd27160}; // indx = 1665
    #10;
    addra = 32'd53312;
    dina = {96'd0, 16'd44252, 16'd39177, 16'd18255, 16'd3539, 16'd12518, 16'd51833, 16'd61756, 16'd57603, 16'd10708, 16'd52926}; // indx = 1666
    #10;
    addra = 32'd53344;
    dina = {96'd0, 16'd33198, 16'd64439, 16'd41258, 16'd4089, 16'd18605, 16'd24475, 16'd20650, 16'd23736, 16'd8451, 16'd44342}; // indx = 1667
    #10;
    addra = 32'd53376;
    dina = {96'd0, 16'd53279, 16'd6882, 16'd11533, 16'd11644, 16'd42452, 16'd62458, 16'd10532, 16'd48832, 16'd51496, 16'd50111}; // indx = 1668
    #10;
    addra = 32'd53408;
    dina = {96'd0, 16'd27777, 16'd33929, 16'd63039, 16'd57221, 16'd11996, 16'd7117, 16'd55804, 16'd65420, 16'd42027, 16'd62652}; // indx = 1669
    #10;
    addra = 32'd53440;
    dina = {96'd0, 16'd51435, 16'd49237, 16'd28203, 16'd19568, 16'd23741, 16'd63628, 16'd40078, 16'd40053, 16'd25776, 16'd53700}; // indx = 1670
    #10;
    addra = 32'd53472;
    dina = {96'd0, 16'd7510, 16'd43188, 16'd3225, 16'd50670, 16'd49422, 16'd22632, 16'd32843, 16'd20695, 16'd54033, 16'd49506}; // indx = 1671
    #10;
    addra = 32'd53504;
    dina = {96'd0, 16'd5076, 16'd30166, 16'd23698, 16'd15070, 16'd27811, 16'd1646, 16'd63992, 16'd48083, 16'd27263, 16'd25935}; // indx = 1672
    #10;
    addra = 32'd53536;
    dina = {96'd0, 16'd29413, 16'd46224, 16'd32403, 16'd46016, 16'd63104, 16'd49995, 16'd3383, 16'd20975, 16'd43608, 16'd59080}; // indx = 1673
    #10;
    addra = 32'd53568;
    dina = {96'd0, 16'd8455, 16'd16542, 16'd59516, 16'd37373, 16'd65343, 16'd16417, 16'd31542, 16'd16408, 16'd41350, 16'd15748}; // indx = 1674
    #10;
    addra = 32'd53600;
    dina = {96'd0, 16'd52776, 16'd49311, 16'd64595, 16'd63376, 16'd28941, 16'd5391, 16'd16270, 16'd4276, 16'd40351, 16'd34488}; // indx = 1675
    #10;
    addra = 32'd53632;
    dina = {96'd0, 16'd40516, 16'd2292, 16'd8049, 16'd42977, 16'd54683, 16'd55507, 16'd23317, 16'd11220, 16'd62404, 16'd10050}; // indx = 1676
    #10;
    addra = 32'd53664;
    dina = {96'd0, 16'd17026, 16'd63417, 16'd57769, 16'd39442, 16'd13482, 16'd54928, 16'd12886, 16'd25043, 16'd9303, 16'd34128}; // indx = 1677
    #10;
    addra = 32'd53696;
    dina = {96'd0, 16'd59824, 16'd37012, 16'd44810, 16'd41541, 16'd21813, 16'd17895, 16'd40000, 16'd52586, 16'd42755, 16'd58537}; // indx = 1678
    #10;
    addra = 32'd53728;
    dina = {96'd0, 16'd42302, 16'd9061, 16'd26196, 16'd26541, 16'd46878, 16'd11989, 16'd16529, 16'd59169, 16'd29265, 16'd45541}; // indx = 1679
    #10;
    addra = 32'd53760;
    dina = {96'd0, 16'd46328, 16'd11470, 16'd57395, 16'd51609, 16'd113, 16'd63045, 16'd28569, 16'd28905, 16'd9565, 16'd21066}; // indx = 1680
    #10;
    addra = 32'd53792;
    dina = {96'd0, 16'd9626, 16'd3289, 16'd8943, 16'd43798, 16'd58495, 16'd57700, 16'd2282, 16'd29334, 16'd24104, 16'd30719}; // indx = 1681
    #10;
    addra = 32'd53824;
    dina = {96'd0, 16'd46162, 16'd49291, 16'd9274, 16'd29649, 16'd7052, 16'd54011, 16'd14695, 16'd26239, 16'd27943, 16'd36426}; // indx = 1682
    #10;
    addra = 32'd53856;
    dina = {96'd0, 16'd2475, 16'd39318, 16'd52126, 16'd53086, 16'd28778, 16'd20960, 16'd5690, 16'd40256, 16'd32776, 16'd32696}; // indx = 1683
    #10;
    addra = 32'd53888;
    dina = {96'd0, 16'd34726, 16'd44388, 16'd3397, 16'd3504, 16'd12851, 16'd25857, 16'd51478, 16'd9377, 16'd32108, 16'd27882}; // indx = 1684
    #10;
    addra = 32'd53920;
    dina = {96'd0, 16'd33571, 16'd14598, 16'd23721, 16'd59166, 16'd23344, 16'd30366, 16'd24016, 16'd34279, 16'd23965, 16'd7215}; // indx = 1685
    #10;
    addra = 32'd53952;
    dina = {96'd0, 16'd63336, 16'd11588, 16'd3726, 16'd62334, 16'd41452, 16'd65511, 16'd61907, 16'd8736, 16'd54627, 16'd1198}; // indx = 1686
    #10;
    addra = 32'd53984;
    dina = {96'd0, 16'd44833, 16'd19806, 16'd12085, 16'd32306, 16'd988, 16'd32759, 16'd63273, 16'd7474, 16'd63175, 16'd2634}; // indx = 1687
    #10;
    addra = 32'd54016;
    dina = {96'd0, 16'd59885, 16'd18124, 16'd24865, 16'd13721, 16'd36172, 16'd25805, 16'd12763, 16'd45777, 16'd28080, 16'd58090}; // indx = 1688
    #10;
    addra = 32'd54048;
    dina = {96'd0, 16'd26293, 16'd48162, 16'd52100, 16'd65143, 16'd56346, 16'd32725, 16'd3369, 16'd21943, 16'd2202, 16'd32019}; // indx = 1689
    #10;
    addra = 32'd54080;
    dina = {96'd0, 16'd32716, 16'd53862, 16'd34915, 16'd54734, 16'd14867, 16'd35581, 16'd22449, 16'd45850, 16'd46816, 16'd20692}; // indx = 1690
    #10;
    addra = 32'd54112;
    dina = {96'd0, 16'd11647, 16'd35811, 16'd50973, 16'd28671, 16'd814, 16'd46216, 16'd46613, 16'd9114, 16'd53026, 16'd38696}; // indx = 1691
    #10;
    addra = 32'd54144;
    dina = {96'd0, 16'd24917, 16'd54348, 16'd5982, 16'd39602, 16'd845, 16'd65184, 16'd5966, 16'd30212, 16'd7807, 16'd60544}; // indx = 1692
    #10;
    addra = 32'd54176;
    dina = {96'd0, 16'd22918, 16'd18919, 16'd18666, 16'd48783, 16'd25195, 16'd38396, 16'd48617, 16'd15596, 16'd15253, 16'd36639}; // indx = 1693
    #10;
    addra = 32'd54208;
    dina = {96'd0, 16'd64743, 16'd31812, 16'd7546, 16'd58473, 16'd4706, 16'd28154, 16'd31722, 16'd29456, 16'd44549, 16'd3777}; // indx = 1694
    #10;
    addra = 32'd54240;
    dina = {96'd0, 16'd40906, 16'd48523, 16'd45122, 16'd14938, 16'd39396, 16'd46123, 16'd39931, 16'd41476, 16'd36018, 16'd51866}; // indx = 1695
    #10;
    addra = 32'd54272;
    dina = {96'd0, 16'd53018, 16'd43024, 16'd26337, 16'd51965, 16'd26878, 16'd40138, 16'd761, 16'd64218, 16'd3624, 16'd21247}; // indx = 1696
    #10;
    addra = 32'd54304;
    dina = {96'd0, 16'd62060, 16'd45885, 16'd62398, 16'd61727, 16'd27571, 16'd51460, 16'd52296, 16'd62273, 16'd20874, 16'd45493}; // indx = 1697
    #10;
    addra = 32'd54336;
    dina = {96'd0, 16'd20679, 16'd20177, 16'd19773, 16'd57958, 16'd20520, 16'd63433, 16'd4075, 16'd11827, 16'd51053, 16'd37552}; // indx = 1698
    #10;
    addra = 32'd54368;
    dina = {96'd0, 16'd3642, 16'd52400, 16'd37234, 16'd29415, 16'd14211, 16'd15045, 16'd404, 16'd22097, 16'd37616, 16'd8622}; // indx = 1699
    #10;
    addra = 32'd54400;
    dina = {96'd0, 16'd56921, 16'd43221, 16'd38959, 16'd31600, 16'd28422, 16'd42878, 16'd50878, 16'd38577, 16'd15614, 16'd31153}; // indx = 1700
    #10;
    addra = 32'd54432;
    dina = {96'd0, 16'd33379, 16'd23454, 16'd46436, 16'd8178, 16'd6468, 16'd43810, 16'd47780, 16'd41979, 16'd56299, 16'd50329}; // indx = 1701
    #10;
    addra = 32'd54464;
    dina = {96'd0, 16'd20568, 16'd25721, 16'd24103, 16'd55956, 16'd62870, 16'd48904, 16'd19677, 16'd19082, 16'd1762, 16'd3344}; // indx = 1702
    #10;
    addra = 32'd54496;
    dina = {96'd0, 16'd23101, 16'd26704, 16'd10898, 16'd37304, 16'd23651, 16'd39817, 16'd56704, 16'd52877, 16'd37572, 16'd54432}; // indx = 1703
    #10;
    addra = 32'd54528;
    dina = {96'd0, 16'd7651, 16'd18089, 16'd38031, 16'd1314, 16'd53734, 16'd12697, 16'd26958, 16'd44142, 16'd31391, 16'd64308}; // indx = 1704
    #10;
    addra = 32'd54560;
    dina = {96'd0, 16'd20848, 16'd13754, 16'd20690, 16'd35961, 16'd41490, 16'd26266, 16'd42133, 16'd19189, 16'd33687, 16'd18842}; // indx = 1705
    #10;
    addra = 32'd54592;
    dina = {96'd0, 16'd59341, 16'd15165, 16'd27247, 16'd4745, 16'd54263, 16'd58362, 16'd51247, 16'd63416, 16'd29773, 16'd34261}; // indx = 1706
    #10;
    addra = 32'd54624;
    dina = {96'd0, 16'd62698, 16'd60510, 16'd43861, 16'd54324, 16'd40825, 16'd29742, 16'd28604, 16'd27584, 16'd61554, 16'd29652}; // indx = 1707
    #10;
    addra = 32'd54656;
    dina = {96'd0, 16'd28116, 16'd57213, 16'd48075, 16'd27814, 16'd42827, 16'd32968, 16'd47023, 16'd5345, 16'd14738, 16'd53649}; // indx = 1708
    #10;
    addra = 32'd54688;
    dina = {96'd0, 16'd21049, 16'd43779, 16'd35828, 16'd52268, 16'd30298, 16'd37785, 16'd15658, 16'd28006, 16'd34024, 16'd53898}; // indx = 1709
    #10;
    addra = 32'd54720;
    dina = {96'd0, 16'd6273, 16'd40093, 16'd29480, 16'd45079, 16'd12946, 16'd15400, 16'd34197, 16'd59625, 16'd44814, 16'd10245}; // indx = 1710
    #10;
    addra = 32'd54752;
    dina = {96'd0, 16'd15715, 16'd61726, 16'd41839, 16'd59141, 16'd55318, 16'd13290, 16'd7098, 16'd65400, 16'd28752, 16'd49204}; // indx = 1711
    #10;
    addra = 32'd54784;
    dina = {96'd0, 16'd3523, 16'd47088, 16'd53594, 16'd53653, 16'd35899, 16'd44853, 16'd5051, 16'd5264, 16'd50374, 16'd38185}; // indx = 1712
    #10;
    addra = 32'd54816;
    dina = {96'd0, 16'd19458, 16'd8636, 16'd65148, 16'd18486, 16'd8403, 16'd16410, 16'd43505, 16'd63109, 16'd65404, 16'd64553}; // indx = 1713
    #10;
    addra = 32'd54848;
    dina = {96'd0, 16'd55783, 16'd56768, 16'd318, 16'd50604, 16'd3016, 16'd30425, 16'd3912, 16'd46443, 16'd8300, 16'd6885}; // indx = 1714
    #10;
    addra = 32'd54880;
    dina = {96'd0, 16'd41461, 16'd54727, 16'd41216, 16'd10212, 16'd16906, 16'd15160, 16'd1706, 16'd32439, 16'd36079, 16'd52411}; // indx = 1715
    #10;
    addra = 32'd54912;
    dina = {96'd0, 16'd46955, 16'd30796, 16'd12555, 16'd17128, 16'd52298, 16'd35031, 16'd14301, 16'd59330, 16'd49573, 16'd37912}; // indx = 1716
    #10;
    addra = 32'd54944;
    dina = {96'd0, 16'd9844, 16'd36375, 16'd64120, 16'd63502, 16'd35175, 16'd3361, 16'd64406, 16'd3864, 16'd42423, 16'd29249}; // indx = 1717
    #10;
    addra = 32'd54976;
    dina = {96'd0, 16'd64893, 16'd28204, 16'd36921, 16'd62198, 16'd28035, 16'd48328, 16'd56062, 16'd17855, 16'd26653, 16'd36856}; // indx = 1718
    #10;
    addra = 32'd55008;
    dina = {96'd0, 16'd13854, 16'd10902, 16'd33928, 16'd64067, 16'd50913, 16'd58177, 16'd22425, 16'd10883, 16'd16811, 16'd50021}; // indx = 1719
    #10;
    addra = 32'd55040;
    dina = {96'd0, 16'd24399, 16'd12695, 16'd10740, 16'd37370, 16'd34106, 16'd3156, 16'd39701, 16'd6204, 16'd24674, 16'd49579}; // indx = 1720
    #10;
    addra = 32'd55072;
    dina = {96'd0, 16'd55822, 16'd41687, 16'd1543, 16'd54798, 16'd32064, 16'd56283, 16'd35716, 16'd16754, 16'd14513, 16'd4872}; // indx = 1721
    #10;
    addra = 32'd55104;
    dina = {96'd0, 16'd25127, 16'd58770, 16'd21654, 16'd49556, 16'd14785, 16'd38742, 16'd13660, 16'd30623, 16'd57090, 16'd28698}; // indx = 1722
    #10;
    addra = 32'd55136;
    dina = {96'd0, 16'd106, 16'd38021, 16'd49257, 16'd47771, 16'd51848, 16'd41009, 16'd2875, 16'd27821, 16'd43739, 16'd54734}; // indx = 1723
    #10;
    addra = 32'd55168;
    dina = {96'd0, 16'd25555, 16'd47776, 16'd27636, 16'd57449, 16'd44029, 16'd33814, 16'd279, 16'd31534, 16'd18603, 16'd51609}; // indx = 1724
    #10;
    addra = 32'd55200;
    dina = {96'd0, 16'd43234, 16'd16641, 16'd20916, 16'd59111, 16'd20055, 16'd32584, 16'd36656, 16'd48744, 16'd39426, 16'd16058}; // indx = 1725
    #10;
    addra = 32'd55232;
    dina = {96'd0, 16'd14179, 16'd37818, 16'd22530, 16'd26403, 16'd39075, 16'd7831, 16'd2560, 16'd60241, 16'd36513, 16'd8526}; // indx = 1726
    #10;
    addra = 32'd55264;
    dina = {96'd0, 16'd59987, 16'd41456, 16'd9462, 16'd50249, 16'd3454, 16'd36372, 16'd37870, 16'd48249, 16'd56915, 16'd6562}; // indx = 1727
    #10;
    addra = 32'd55296;
    dina = {96'd0, 16'd4125, 16'd14507, 16'd58544, 16'd36601, 16'd60560, 16'd55617, 16'd32458, 16'd3039, 16'd57048, 16'd13614}; // indx = 1728
    #10;
    addra = 32'd55328;
    dina = {96'd0, 16'd37150, 16'd37390, 16'd39142, 16'd43036, 16'd5935, 16'd31857, 16'd52457, 16'd15740, 16'd32802, 16'd54364}; // indx = 1729
    #10;
    addra = 32'd55360;
    dina = {96'd0, 16'd39429, 16'd20991, 16'd17642, 16'd58101, 16'd57391, 16'd43265, 16'd35026, 16'd8930, 16'd13665, 16'd55030}; // indx = 1730
    #10;
    addra = 32'd55392;
    dina = {96'd0, 16'd64118, 16'd35938, 16'd21350, 16'd9001, 16'd49163, 16'd50297, 16'd22809, 16'd14620, 16'd34383, 16'd41105}; // indx = 1731
    #10;
    addra = 32'd55424;
    dina = {96'd0, 16'd42488, 16'd44133, 16'd43528, 16'd1295, 16'd19992, 16'd44653, 16'd1548, 16'd49451, 16'd61991, 16'd41843}; // indx = 1732
    #10;
    addra = 32'd55456;
    dina = {96'd0, 16'd52392, 16'd62215, 16'd23037, 16'd7689, 16'd17182, 16'd46237, 16'd46416, 16'd46185, 16'd35715, 16'd40786}; // indx = 1733
    #10;
    addra = 32'd55488;
    dina = {96'd0, 16'd15604, 16'd21862, 16'd43440, 16'd34063, 16'd14390, 16'd3435, 16'd50191, 16'd20101, 16'd45070, 16'd23196}; // indx = 1734
    #10;
    addra = 32'd55520;
    dina = {96'd0, 16'd36651, 16'd40262, 16'd23751, 16'd35798, 16'd52238, 16'd54889, 16'd43169, 16'd63666, 16'd26634, 16'd59934}; // indx = 1735
    #10;
    addra = 32'd55552;
    dina = {96'd0, 16'd34067, 16'd36419, 16'd49519, 16'd42247, 16'd44728, 16'd57312, 16'd22989, 16'd61457, 16'd62774, 16'd14897}; // indx = 1736
    #10;
    addra = 32'd55584;
    dina = {96'd0, 16'd3764, 16'd49198, 16'd7113, 16'd48283, 16'd6858, 16'd32973, 16'd54747, 16'd59618, 16'd62809, 16'd10621}; // indx = 1737
    #10;
    addra = 32'd55616;
    dina = {96'd0, 16'd25, 16'd48807, 16'd20386, 16'd36502, 16'd36281, 16'd46063, 16'd48685, 16'd11115, 16'd33897, 16'd62529}; // indx = 1738
    #10;
    addra = 32'd55648;
    dina = {96'd0, 16'd45611, 16'd54014, 16'd48832, 16'd49007, 16'd58117, 16'd52964, 16'd694, 16'd37366, 16'd19690, 16'd62074}; // indx = 1739
    #10;
    addra = 32'd55680;
    dina = {96'd0, 16'd13982, 16'd40691, 16'd6609, 16'd28703, 16'd38182, 16'd21117, 16'd2474, 16'd58175, 16'd60672, 16'd1717}; // indx = 1740
    #10;
    addra = 32'd55712;
    dina = {96'd0, 16'd22356, 16'd48745, 16'd55523, 16'd36701, 16'd64186, 16'd22771, 16'd51976, 16'd44585, 16'd42408, 16'd57265}; // indx = 1741
    #10;
    addra = 32'd55744;
    dina = {96'd0, 16'd17024, 16'd37059, 16'd18504, 16'd35552, 16'd45931, 16'd39721, 16'd56348, 16'd62330, 16'd10520, 16'd44453}; // indx = 1742
    #10;
    addra = 32'd55776;
    dina = {96'd0, 16'd32847, 16'd64886, 16'd4759, 16'd29649, 16'd15326, 16'd42432, 16'd35825, 16'd10002, 16'd33579, 16'd54251}; // indx = 1743
    #10;
    addra = 32'd55808;
    dina = {96'd0, 16'd12050, 16'd38190, 16'd46006, 16'd14502, 16'd5730, 16'd25112, 16'd19486, 16'd44433, 16'd18051, 16'd1346}; // indx = 1744
    #10;
    addra = 32'd55840;
    dina = {96'd0, 16'd38771, 16'd15561, 16'd19164, 16'd29717, 16'd22758, 16'd48037, 16'd6544, 16'd24826, 16'd63933, 16'd22459}; // indx = 1745
    #10;
    addra = 32'd55872;
    dina = {96'd0, 16'd23563, 16'd34233, 16'd7478, 16'd49531, 16'd44955, 16'd1398, 16'd54326, 16'd60932, 16'd27254, 16'd51512}; // indx = 1746
    #10;
    addra = 32'd55904;
    dina = {96'd0, 16'd27773, 16'd38860, 16'd14952, 16'd6527, 16'd8473, 16'd40575, 16'd16225, 16'd32156, 16'd5940, 16'd49954}; // indx = 1747
    #10;
    addra = 32'd55936;
    dina = {96'd0, 16'd63883, 16'd10162, 16'd30440, 16'd21926, 16'd40434, 16'd9867, 16'd29284, 16'd13949, 16'd464, 16'd32695}; // indx = 1748
    #10;
    addra = 32'd55968;
    dina = {96'd0, 16'd6631, 16'd21625, 16'd34960, 16'd40904, 16'd392, 16'd32621, 16'd34605, 16'd40109, 16'd3379, 16'd45093}; // indx = 1749
    #10;
    addra = 32'd56000;
    dina = {96'd0, 16'd52588, 16'd45534, 16'd54150, 16'd51265, 16'd45627, 16'd15355, 16'd27618, 16'd8542, 16'd17549, 16'd56771}; // indx = 1750
    #10;
    addra = 32'd56032;
    dina = {96'd0, 16'd43066, 16'd58321, 16'd10722, 16'd31997, 16'd18482, 16'd24190, 16'd26083, 16'd48835, 16'd9041, 16'd40520}; // indx = 1751
    #10;
    addra = 32'd56064;
    dina = {96'd0, 16'd44488, 16'd45762, 16'd53114, 16'd34965, 16'd29688, 16'd56029, 16'd1749, 16'd4349, 16'd60746, 16'd29982}; // indx = 1752
    #10;
    addra = 32'd56096;
    dina = {96'd0, 16'd24312, 16'd58328, 16'd12239, 16'd27489, 16'd32702, 16'd3235, 16'd359, 16'd61782, 16'd3987, 16'd11701}; // indx = 1753
    #10;
    addra = 32'd56128;
    dina = {96'd0, 16'd3258, 16'd61842, 16'd44337, 16'd18478, 16'd17241, 16'd2100, 16'd16214, 16'd37773, 16'd24792, 16'd2542}; // indx = 1754
    #10;
    addra = 32'd56160;
    dina = {96'd0, 16'd34352, 16'd30091, 16'd55258, 16'd21974, 16'd32155, 16'd11500, 16'd15942, 16'd19810, 16'd16284, 16'd47780}; // indx = 1755
    #10;
    addra = 32'd56192;
    dina = {96'd0, 16'd7524, 16'd31211, 16'd15759, 16'd32960, 16'd29811, 16'd59043, 16'd12890, 16'd11653, 16'd63752, 16'd3851}; // indx = 1756
    #10;
    addra = 32'd56224;
    dina = {96'd0, 16'd45910, 16'd18996, 16'd11645, 16'd31287, 16'd48499, 16'd43361, 16'd48591, 16'd29471, 16'd29953, 16'd53309}; // indx = 1757
    #10;
    addra = 32'd56256;
    dina = {96'd0, 16'd37417, 16'd28484, 16'd27458, 16'd23056, 16'd33136, 16'd44882, 16'd60499, 16'd41862, 16'd3272, 16'd30485}; // indx = 1758
    #10;
    addra = 32'd56288;
    dina = {96'd0, 16'd23544, 16'd53229, 16'd579, 16'd36013, 16'd62857, 16'd19341, 16'd65468, 16'd65018, 16'd23059, 16'd19893}; // indx = 1759
    #10;
    addra = 32'd56320;
    dina = {96'd0, 16'd24612, 16'd53306, 16'd46064, 16'd39122, 16'd27615, 16'd57524, 16'd59428, 16'd47259, 16'd32108, 16'd51162}; // indx = 1760
    #10;
    addra = 32'd56352;
    dina = {96'd0, 16'd32012, 16'd14171, 16'd9904, 16'd19611, 16'd26897, 16'd22111, 16'd41384, 16'd43382, 16'd24424, 16'd57097}; // indx = 1761
    #10;
    addra = 32'd56384;
    dina = {96'd0, 16'd36887, 16'd23097, 16'd9611, 16'd15060, 16'd55150, 16'd30375, 16'd30348, 16'd18056, 16'd8023, 16'd7565}; // indx = 1762
    #10;
    addra = 32'd56416;
    dina = {96'd0, 16'd9506, 16'd14331, 16'd21197, 16'd22414, 16'd54542, 16'd250, 16'd22170, 16'd23034, 16'd14257, 16'd24005}; // indx = 1763
    #10;
    addra = 32'd56448;
    dina = {96'd0, 16'd61081, 16'd23025, 16'd21496, 16'd32453, 16'd7860, 16'd8490, 16'd18522, 16'd62960, 16'd12424, 16'd3840}; // indx = 1764
    #10;
    addra = 32'd56480;
    dina = {96'd0, 16'd1289, 16'd11084, 16'd10811, 16'd13839, 16'd38825, 16'd19065, 16'd55961, 16'd12602, 16'd34784, 16'd23879}; // indx = 1765
    #10;
    addra = 32'd56512;
    dina = {96'd0, 16'd57820, 16'd25195, 16'd49554, 16'd24291, 16'd29360, 16'd52992, 16'd56419, 16'd11178, 16'd15490, 16'd9495}; // indx = 1766
    #10;
    addra = 32'd56544;
    dina = {96'd0, 16'd16572, 16'd30456, 16'd21766, 16'd55617, 16'd58627, 16'd2125, 16'd34193, 16'd764, 16'd60137, 16'd42932}; // indx = 1767
    #10;
    addra = 32'd56576;
    dina = {96'd0, 16'd38317, 16'd63314, 16'd39266, 16'd20904, 16'd48348, 16'd36228, 16'd36967, 16'd36275, 16'd28997, 16'd13196}; // indx = 1768
    #10;
    addra = 32'd56608;
    dina = {96'd0, 16'd55825, 16'd13943, 16'd33651, 16'd41707, 16'd61132, 16'd15112, 16'd34481, 16'd19672, 16'd103, 16'd3897}; // indx = 1769
    #10;
    addra = 32'd56640;
    dina = {96'd0, 16'd34502, 16'd39624, 16'd63183, 16'd28510, 16'd57053, 16'd19399, 16'd59214, 16'd11241, 16'd22944, 16'd9310}; // indx = 1770
    #10;
    addra = 32'd56672;
    dina = {96'd0, 16'd64473, 16'd32775, 16'd32104, 16'd56996, 16'd5159, 16'd31038, 16'd40189, 16'd12194, 16'd26730, 16'd33682}; // indx = 1771
    #10;
    addra = 32'd56704;
    dina = {96'd0, 16'd47373, 16'd8727, 16'd38125, 16'd51288, 16'd55695, 16'd27100, 16'd21478, 16'd18672, 16'd4739, 16'd20140}; // indx = 1772
    #10;
    addra = 32'd56736;
    dina = {96'd0, 16'd56322, 16'd18399, 16'd39328, 16'd65232, 16'd6355, 16'd471, 16'd56236, 16'd48098, 16'd14556, 16'd687}; // indx = 1773
    #10;
    addra = 32'd56768;
    dina = {96'd0, 16'd35556, 16'd27016, 16'd17197, 16'd60072, 16'd52404, 16'd54687, 16'd12487, 16'd53192, 16'd24459, 16'd52529}; // indx = 1774
    #10;
    addra = 32'd56800;
    dina = {96'd0, 16'd53074, 16'd19760, 16'd59865, 16'd65459, 16'd36099, 16'd33949, 16'd56704, 16'd9515, 16'd27276, 16'd64681}; // indx = 1775
    #10;
    addra = 32'd56832;
    dina = {96'd0, 16'd44187, 16'd42527, 16'd34105, 16'd19573, 16'd49326, 16'd60969, 16'd42678, 16'd11427, 16'd34667, 16'd22819}; // indx = 1776
    #10;
    addra = 32'd56864;
    dina = {96'd0, 16'd43993, 16'd40167, 16'd1391, 16'd59950, 16'd4249, 16'd48024, 16'd9639, 16'd59351, 16'd8917, 16'd2675}; // indx = 1777
    #10;
    addra = 32'd56896;
    dina = {96'd0, 16'd335, 16'd61046, 16'd37670, 16'd31845, 16'd49170, 16'd11509, 16'd33881, 16'd32116, 16'd4925, 16'd2053}; // indx = 1778
    #10;
    addra = 32'd56928;
    dina = {96'd0, 16'd35973, 16'd45150, 16'd57235, 16'd16100, 16'd62350, 16'd44404, 16'd7899, 16'd28328, 16'd10326, 16'd35061}; // indx = 1779
    #10;
    addra = 32'd56960;
    dina = {96'd0, 16'd33201, 16'd48615, 16'd29299, 16'd41703, 16'd58641, 16'd57810, 16'd49998, 16'd7723, 16'd55099, 16'd61801}; // indx = 1780
    #10;
    addra = 32'd56992;
    dina = {96'd0, 16'd18234, 16'd39448, 16'd58590, 16'd63870, 16'd18329, 16'd2339, 16'd10937, 16'd26313, 16'd49413, 16'd36771}; // indx = 1781
    #10;
    addra = 32'd57024;
    dina = {96'd0, 16'd17377, 16'd44946, 16'd22304, 16'd7060, 16'd33891, 16'd17853, 16'd34345, 16'd18519, 16'd25762, 16'd31860}; // indx = 1782
    #10;
    addra = 32'd57056;
    dina = {96'd0, 16'd14639, 16'd46995, 16'd11076, 16'd26752, 16'd2135, 16'd54199, 16'd53518, 16'd52333, 16'd5175, 16'd49425}; // indx = 1783
    #10;
    addra = 32'd57088;
    dina = {96'd0, 16'd4355, 16'd17082, 16'd20735, 16'd24562, 16'd8968, 16'd30199, 16'd45253, 16'd41429, 16'd6614, 16'd3134}; // indx = 1784
    #10;
    addra = 32'd57120;
    dina = {96'd0, 16'd9914, 16'd38606, 16'd46343, 16'd7094, 16'd50806, 16'd50335, 16'd8931, 16'd11604, 16'd63493, 16'd56922}; // indx = 1785
    #10;
    addra = 32'd57152;
    dina = {96'd0, 16'd7140, 16'd52310, 16'd28248, 16'd50049, 16'd33035, 16'd23240, 16'd65273, 16'd39613, 16'd6469, 16'd21905}; // indx = 1786
    #10;
    addra = 32'd57184;
    dina = {96'd0, 16'd59319, 16'd41719, 16'd52808, 16'd11477, 16'd41637, 16'd22156, 16'd29318, 16'd17212, 16'd62658, 16'd29291}; // indx = 1787
    #10;
    addra = 32'd57216;
    dina = {96'd0, 16'd364, 16'd64257, 16'd36818, 16'd41822, 16'd22097, 16'd30706, 16'd18539, 16'd24797, 16'd58267, 16'd24778}; // indx = 1788
    #10;
    addra = 32'd57248;
    dina = {96'd0, 16'd62308, 16'd46397, 16'd61782, 16'd35439, 16'd27234, 16'd28704, 16'd54589, 16'd54271, 16'd62978, 16'd36559}; // indx = 1789
    #10;
    addra = 32'd57280;
    dina = {96'd0, 16'd50652, 16'd417, 16'd53289, 16'd12097, 16'd33589, 16'd43680, 16'd19916, 16'd15417, 16'd60187, 16'd51223}; // indx = 1790
    #10;
    addra = 32'd57312;
    dina = {96'd0, 16'd3136, 16'd39358, 16'd32967, 16'd30973, 16'd33830, 16'd39634, 16'd11249, 16'd1285, 16'd4311, 16'd36684}; // indx = 1791
    #10;
    addra = 32'd57344;
    dina = {96'd0, 16'd56801, 16'd55819, 16'd11513, 16'd30109, 16'd27862, 16'd53099, 16'd31127, 16'd12778, 16'd47478, 16'd12898}; // indx = 1792
    #10;
    addra = 32'd57376;
    dina = {96'd0, 16'd50811, 16'd40682, 16'd63606, 16'd29452, 16'd30151, 16'd4581, 16'd8299, 16'd34071, 16'd53619, 16'd30186}; // indx = 1793
    #10;
    addra = 32'd57408;
    dina = {96'd0, 16'd35418, 16'd22305, 16'd47905, 16'd64459, 16'd53163, 16'd20674, 16'd17090, 16'd5994, 16'd28765, 16'd21853}; // indx = 1794
    #10;
    addra = 32'd57440;
    dina = {96'd0, 16'd27417, 16'd61816, 16'd20019, 16'd19474, 16'd58541, 16'd13265, 16'd1396, 16'd21692, 16'd10813, 16'd60131}; // indx = 1795
    #10;
    addra = 32'd57472;
    dina = {96'd0, 16'd40199, 16'd33971, 16'd24861, 16'd44536, 16'd29721, 16'd19314, 16'd12812, 16'd20510, 16'd54284, 16'd25312}; // indx = 1796
    #10;
    addra = 32'd57504;
    dina = {96'd0, 16'd8833, 16'd53692, 16'd31067, 16'd26167, 16'd54818, 16'd44762, 16'd28352, 16'd49564, 16'd34756, 16'd13762}; // indx = 1797
    #10;
    addra = 32'd57536;
    dina = {96'd0, 16'd50379, 16'd50137, 16'd16783, 16'd38005, 16'd25446, 16'd15805, 16'd11579, 16'd51105, 16'd56637, 16'd21793}; // indx = 1798
    #10;
    addra = 32'd57568;
    dina = {96'd0, 16'd61913, 16'd44148, 16'd63672, 16'd54017, 16'd14910, 16'd24265, 16'd6375, 16'd32386, 16'd49783, 16'd8319}; // indx = 1799
    #10;
    addra = 32'd57600;
    dina = {96'd0, 16'd44772, 16'd8045, 16'd3688, 16'd55059, 16'd18102, 16'd29652, 16'd8689, 16'd55672, 16'd25759, 16'd12825}; // indx = 1800
    #10;
    addra = 32'd57632;
    dina = {96'd0, 16'd26827, 16'd7680, 16'd40553, 16'd32012, 16'd37411, 16'd21520, 16'd38365, 16'd35985, 16'd48719, 16'd18512}; // indx = 1801
    #10;
    addra = 32'd57664;
    dina = {96'd0, 16'd29164, 16'd46986, 16'd42235, 16'd23451, 16'd38354, 16'd9751, 16'd23125, 16'd75, 16'd56056, 16'd27645}; // indx = 1802
    #10;
    addra = 32'd57696;
    dina = {96'd0, 16'd1770, 16'd61255, 16'd49921, 16'd59683, 16'd65024, 16'd62819, 16'd6993, 16'd65209, 16'd16523, 16'd49389}; // indx = 1803
    #10;
    addra = 32'd57728;
    dina = {96'd0, 16'd27533, 16'd25052, 16'd12634, 16'd26776, 16'd20797, 16'd33524, 16'd18885, 16'd39248, 16'd60397, 16'd24307}; // indx = 1804
    #10;
    addra = 32'd57760;
    dina = {96'd0, 16'd47687, 16'd47860, 16'd9491, 16'd11832, 16'd14732, 16'd38155, 16'd23582, 16'd42857, 16'd46015, 16'd36638}; // indx = 1805
    #10;
    addra = 32'd57792;
    dina = {96'd0, 16'd50293, 16'd48578, 16'd15545, 16'd64225, 16'd54086, 16'd50366, 16'd34269, 16'd24151, 16'd26397, 16'd31525}; // indx = 1806
    #10;
    addra = 32'd57824;
    dina = {96'd0, 16'd19590, 16'd22916, 16'd36636, 16'd39705, 16'd47047, 16'd35283, 16'd53372, 16'd64337, 16'd45557, 16'd22121}; // indx = 1807
    #10;
    addra = 32'd57856;
    dina = {96'd0, 16'd42566, 16'd55995, 16'd24127, 16'd48694, 16'd11419, 16'd39452, 16'd56238, 16'd38633, 16'd10231, 16'd49112}; // indx = 1808
    #10;
    addra = 32'd57888;
    dina = {96'd0, 16'd19123, 16'd19472, 16'd57506, 16'd6704, 16'd45449, 16'd12677, 16'd36680, 16'd11301, 16'd1300, 16'd51022}; // indx = 1809
    #10;
    addra = 32'd57920;
    dina = {96'd0, 16'd38651, 16'd46854, 16'd56256, 16'd19812, 16'd12380, 16'd44094, 16'd42658, 16'd25606, 16'd32702, 16'd52492}; // indx = 1810
    #10;
    addra = 32'd57952;
    dina = {96'd0, 16'd9051, 16'd16899, 16'd50196, 16'd11057, 16'd65043, 16'd43728, 16'd9161, 16'd44941, 16'd40783, 16'd9828}; // indx = 1811
    #10;
    addra = 32'd57984;
    dina = {96'd0, 16'd9427, 16'd62787, 16'd56119, 16'd41113, 16'd32355, 16'd41837, 16'd2972, 16'd26399, 16'd54298, 16'd57493}; // indx = 1812
    #10;
    addra = 32'd58016;
    dina = {96'd0, 16'd22847, 16'd25915, 16'd64710, 16'd53909, 16'd61964, 16'd19575, 16'd23535, 16'd8107, 16'd9854, 16'd64867}; // indx = 1813
    #10;
    addra = 32'd58048;
    dina = {96'd0, 16'd28276, 16'd60153, 16'd46028, 16'd5927, 16'd62795, 16'd39425, 16'd55635, 16'd30735, 16'd46594, 16'd57365}; // indx = 1814
    #10;
    addra = 32'd58080;
    dina = {96'd0, 16'd56319, 16'd20082, 16'd54120, 16'd41148, 16'd27253, 16'd62978, 16'd22131, 16'd8729, 16'd20062, 16'd6888}; // indx = 1815
    #10;
    addra = 32'd58112;
    dina = {96'd0, 16'd40935, 16'd47947, 16'd6555, 16'd5172, 16'd53530, 16'd18177, 16'd33217, 16'd52908, 16'd16388, 16'd60150}; // indx = 1816
    #10;
    addra = 32'd58144;
    dina = {96'd0, 16'd2293, 16'd36344, 16'd2574, 16'd15282, 16'd34590, 16'd9221, 16'd47766, 16'd15503, 16'd41838, 16'd48671}; // indx = 1817
    #10;
    addra = 32'd58176;
    dina = {96'd0, 16'd65375, 16'd37767, 16'd40822, 16'd21073, 16'd27878, 16'd62742, 16'd19256, 16'd30881, 16'd28830, 16'd3601}; // indx = 1818
    #10;
    addra = 32'd58208;
    dina = {96'd0, 16'd24057, 16'd31300, 16'd42694, 16'd5854, 16'd1907, 16'd42625, 16'd6300, 16'd42790, 16'd40688, 16'd34256}; // indx = 1819
    #10;
    addra = 32'd58240;
    dina = {96'd0, 16'd41591, 16'd7381, 16'd33759, 16'd15464, 16'd33742, 16'd18661, 16'd33377, 16'd61365, 16'd36758, 16'd11092}; // indx = 1820
    #10;
    addra = 32'd58272;
    dina = {96'd0, 16'd8096, 16'd63362, 16'd28485, 16'd16938, 16'd1054, 16'd32439, 16'd4630, 16'd7105, 16'd24054, 16'd64194}; // indx = 1821
    #10;
    addra = 32'd58304;
    dina = {96'd0, 16'd22274, 16'd55057, 16'd29793, 16'd57640, 16'd33778, 16'd60901, 16'd26586, 16'd58372, 16'd10217, 16'd7276}; // indx = 1822
    #10;
    addra = 32'd58336;
    dina = {96'd0, 16'd57758, 16'd50235, 16'd63916, 16'd65295, 16'd9292, 16'd64279, 16'd41882, 16'd46114, 16'd1854, 16'd32619}; // indx = 1823
    #10;
    addra = 32'd58368;
    dina = {96'd0, 16'd34583, 16'd719, 16'd9528, 16'd31515, 16'd35426, 16'd51129, 16'd61947, 16'd8406, 16'd59557, 16'd50514}; // indx = 1824
    #10;
    addra = 32'd58400;
    dina = {96'd0, 16'd7665, 16'd47859, 16'd4971, 16'd17540, 16'd17460, 16'd43790, 16'd48994, 16'd57072, 16'd5594, 16'd22217}; // indx = 1825
    #10;
    addra = 32'd58432;
    dina = {96'd0, 16'd29183, 16'd63205, 16'd64060, 16'd52385, 16'd24095, 16'd50567, 16'd39819, 16'd5222, 16'd16141, 16'd13128}; // indx = 1826
    #10;
    addra = 32'd58464;
    dina = {96'd0, 16'd14647, 16'd54640, 16'd22696, 16'd41168, 16'd2929, 16'd15007, 16'd15720, 16'd33908, 16'd29296, 16'd2268}; // indx = 1827
    #10;
    addra = 32'd58496;
    dina = {96'd0, 16'd56134, 16'd21484, 16'd3738, 16'd31051, 16'd1747, 16'd53833, 16'd1699, 16'd20446, 16'd5340, 16'd2644}; // indx = 1828
    #10;
    addra = 32'd58528;
    dina = {96'd0, 16'd20526, 16'd23783, 16'd64215, 16'd45, 16'd62806, 16'd23889, 16'd59661, 16'd23726, 16'd55500, 16'd61383}; // indx = 1829
    #10;
    addra = 32'd58560;
    dina = {96'd0, 16'd45713, 16'd12324, 16'd9591, 16'd48741, 16'd31772, 16'd20289, 16'd18764, 16'd41906, 16'd19441, 16'd26069}; // indx = 1830
    #10;
    addra = 32'd58592;
    dina = {96'd0, 16'd13606, 16'd34344, 16'd894, 16'd44946, 16'd18212, 16'd33635, 16'd30435, 16'd30262, 16'd49550, 16'd14114}; // indx = 1831
    #10;
    addra = 32'd58624;
    dina = {96'd0, 16'd57167, 16'd8355, 16'd55925, 16'd9074, 16'd15302, 16'd41734, 16'd56190, 16'd51313, 16'd40324, 16'd5090}; // indx = 1832
    #10;
    addra = 32'd58656;
    dina = {96'd0, 16'd53537, 16'd49176, 16'd53688, 16'd16444, 16'd38428, 16'd64504, 16'd33836, 16'd6834, 16'd29827, 16'd33987}; // indx = 1833
    #10;
    addra = 32'd58688;
    dina = {96'd0, 16'd57544, 16'd12559, 16'd3208, 16'd35720, 16'd37096, 16'd54415, 16'd9775, 16'd46017, 16'd45571, 16'd43702}; // indx = 1834
    #10;
    addra = 32'd58720;
    dina = {96'd0, 16'd46222, 16'd13428, 16'd24871, 16'd25847, 16'd30518, 16'd57598, 16'd15573, 16'd53938, 16'd48472, 16'd8090}; // indx = 1835
    #10;
    addra = 32'd58752;
    dina = {96'd0, 16'd37352, 16'd34818, 16'd8775, 16'd54512, 16'd7434, 16'd16995, 16'd28929, 16'd54535, 16'd39874, 16'd47150}; // indx = 1836
    #10;
    addra = 32'd58784;
    dina = {96'd0, 16'd2719, 16'd32968, 16'd55809, 16'd52143, 16'd9259, 16'd65433, 16'd22598, 16'd14299, 16'd46097, 16'd53765}; // indx = 1837
    #10;
    addra = 32'd58816;
    dina = {96'd0, 16'd38044, 16'd37605, 16'd62077, 16'd44294, 16'd7765, 16'd45250, 16'd52299, 16'd9332, 16'd55281, 16'd56452}; // indx = 1838
    #10;
    addra = 32'd58848;
    dina = {96'd0, 16'd14849, 16'd45085, 16'd21427, 16'd8756, 16'd6667, 16'd4136, 16'd13751, 16'd32529, 16'd23458, 16'd41361}; // indx = 1839
    #10;
    addra = 32'd58880;
    dina = {96'd0, 16'd50348, 16'd59287, 16'd43421, 16'd55753, 16'd57286, 16'd39109, 16'd47575, 16'd24322, 16'd13168, 16'd5880}; // indx = 1840
    #10;
    addra = 32'd58912;
    dina = {96'd0, 16'd42392, 16'd30358, 16'd12951, 16'd33815, 16'd64773, 16'd56244, 16'd16479, 16'd24384, 16'd53478, 16'd4918}; // indx = 1841
    #10;
    addra = 32'd58944;
    dina = {96'd0, 16'd19902, 16'd64230, 16'd7702, 16'd45081, 16'd54558, 16'd32806, 16'd55954, 16'd48002, 16'd64621, 16'd15907}; // indx = 1842
    #10;
    addra = 32'd58976;
    dina = {96'd0, 16'd59020, 16'd37912, 16'd64416, 16'd24888, 16'd3286, 16'd51240, 16'd58042, 16'd27157, 16'd31098, 16'd45655}; // indx = 1843
    #10;
    addra = 32'd59008;
    dina = {96'd0, 16'd59381, 16'd25751, 16'd30951, 16'd19789, 16'd16908, 16'd63588, 16'd41358, 16'd54040, 16'd32616, 16'd6405}; // indx = 1844
    #10;
    addra = 32'd59040;
    dina = {96'd0, 16'd12532, 16'd63736, 16'd38381, 16'd21530, 16'd31008, 16'd31208, 16'd15738, 16'd2060, 16'd410, 16'd41346}; // indx = 1845
    #10;
    addra = 32'd59072;
    dina = {96'd0, 16'd57350, 16'd24146, 16'd13755, 16'd42955, 16'd30756, 16'd62075, 16'd39666, 16'd18471, 16'd45048, 16'd44573}; // indx = 1846
    #10;
    addra = 32'd59104;
    dina = {96'd0, 16'd60325, 16'd45283, 16'd64509, 16'd64495, 16'd55763, 16'd2350, 16'd26174, 16'd62838, 16'd16133, 16'd30079}; // indx = 1847
    #10;
    addra = 32'd59136;
    dina = {96'd0, 16'd64798, 16'd10337, 16'd19188, 16'd10662, 16'd39636, 16'd21142, 16'd11366, 16'd14249, 16'd58932, 16'd24928}; // indx = 1848
    #10;
    addra = 32'd59168;
    dina = {96'd0, 16'd53045, 16'd50987, 16'd23277, 16'd25342, 16'd13915, 16'd63904, 16'd57939, 16'd10957, 16'd46445, 16'd17228}; // indx = 1849
    #10;
    addra = 32'd59200;
    dina = {96'd0, 16'd64954, 16'd64804, 16'd48476, 16'd4560, 16'd2761, 16'd21219, 16'd1597, 16'd43882, 16'd13295, 16'd38543}; // indx = 1850
    #10;
    addra = 32'd59232;
    dina = {96'd0, 16'd27664, 16'd24760, 16'd10717, 16'd4027, 16'd22053, 16'd42104, 16'd60847, 16'd21387, 16'd11507, 16'd36435}; // indx = 1851
    #10;
    addra = 32'd59264;
    dina = {96'd0, 16'd26088, 16'd57009, 16'd63745, 16'd46874, 16'd28794, 16'd3749, 16'd10756, 16'd24018, 16'd64039, 16'd37014}; // indx = 1852
    #10;
    addra = 32'd59296;
    dina = {96'd0, 16'd36082, 16'd48702, 16'd49457, 16'd28383, 16'd8247, 16'd64644, 16'd5610, 16'd6177, 16'd19152, 16'd36094}; // indx = 1853
    #10;
    addra = 32'd59328;
    dina = {96'd0, 16'd34163, 16'd10134, 16'd21774, 16'd2708, 16'd32805, 16'd15418, 16'd21041, 16'd60828, 16'd12143, 16'd53842}; // indx = 1854
    #10;
    addra = 32'd59360;
    dina = {96'd0, 16'd12179, 16'd42741, 16'd15118, 16'd5967, 16'd25210, 16'd50234, 16'd38977, 16'd57584, 16'd28537, 16'd42142}; // indx = 1855
    #10;
    addra = 32'd59392;
    dina = {96'd0, 16'd22098, 16'd11588, 16'd37197, 16'd6919, 16'd21114, 16'd32584, 16'd32507, 16'd32201, 16'd43727, 16'd2785}; // indx = 1856
    #10;
    addra = 32'd59424;
    dina = {96'd0, 16'd29271, 16'd45760, 16'd42958, 16'd23563, 16'd47515, 16'd22955, 16'd15455, 16'd35492, 16'd4677, 16'd50882}; // indx = 1857
    #10;
    addra = 32'd59456;
    dina = {96'd0, 16'd42114, 16'd42964, 16'd44806, 16'd54685, 16'd1773, 16'd56849, 16'd23396, 16'd61341, 16'd22147, 16'd38403}; // indx = 1858
    #10;
    addra = 32'd59488;
    dina = {96'd0, 16'd17281, 16'd28228, 16'd5409, 16'd63057, 16'd35289, 16'd2537, 16'd26616, 16'd9065, 16'd52517, 16'd9924}; // indx = 1859
    #10;
    addra = 32'd59520;
    dina = {96'd0, 16'd60748, 16'd14011, 16'd35390, 16'd5176, 16'd19580, 16'd39121, 16'd60453, 16'd23874, 16'd11267, 16'd64517}; // indx = 1860
    #10;
    addra = 32'd59552;
    dina = {96'd0, 16'd28335, 16'd60382, 16'd52018, 16'd37031, 16'd53522, 16'd40066, 16'd54423, 16'd7883, 16'd428, 16'd58324}; // indx = 1861
    #10;
    addra = 32'd59584;
    dina = {96'd0, 16'd9454, 16'd34501, 16'd45954, 16'd1301, 16'd5920, 16'd14532, 16'd47933, 16'd60046, 16'd26703, 16'd54744}; // indx = 1862
    #10;
    addra = 32'd59616;
    dina = {96'd0, 16'd1952, 16'd37688, 16'd46093, 16'd29926, 16'd57547, 16'd16911, 16'd6038, 16'd31248, 16'd14869, 16'd32977}; // indx = 1863
    #10;
    addra = 32'd59648;
    dina = {96'd0, 16'd7541, 16'd24073, 16'd35579, 16'd9859, 16'd21724, 16'd6272, 16'd4790, 16'd44053, 16'd35153, 16'd135}; // indx = 1864
    #10;
    addra = 32'd59680;
    dina = {96'd0, 16'd55559, 16'd13545, 16'd11280, 16'd25643, 16'd52882, 16'd21442, 16'd17531, 16'd22894, 16'd6572, 16'd34726}; // indx = 1865
    #10;
    addra = 32'd59712;
    dina = {96'd0, 16'd28809, 16'd63091, 16'd41444, 16'd31078, 16'd50455, 16'd19279, 16'd25220, 16'd57240, 16'd27961, 16'd57446}; // indx = 1866
    #10;
    addra = 32'd59744;
    dina = {96'd0, 16'd39814, 16'd2537, 16'd22704, 16'd29555, 16'd62412, 16'd47788, 16'd29405, 16'd47150, 16'd19534, 16'd6019}; // indx = 1867
    #10;
    addra = 32'd59776;
    dina = {96'd0, 16'd52141, 16'd17509, 16'd15539, 16'd64829, 16'd25539, 16'd52052, 16'd1400, 16'd25865, 16'd29711, 16'd18871}; // indx = 1868
    #10;
    addra = 32'd59808;
    dina = {96'd0, 16'd44897, 16'd3539, 16'd57312, 16'd47636, 16'd37115, 16'd45790, 16'd2935, 16'd43321, 16'd35556, 16'd54073}; // indx = 1869
    #10;
    addra = 32'd59840;
    dina = {96'd0, 16'd31223, 16'd19031, 16'd57696, 16'd52861, 16'd22266, 16'd62503, 16'd8651, 16'd28632, 16'd18896, 16'd52657}; // indx = 1870
    #10;
    addra = 32'd59872;
    dina = {96'd0, 16'd47102, 16'd28600, 16'd55183, 16'd47144, 16'd572, 16'd59406, 16'd50787, 16'd51210, 16'd59679, 16'd1130}; // indx = 1871
    #10;
    addra = 32'd59904;
    dina = {96'd0, 16'd63208, 16'd241, 16'd6366, 16'd47901, 16'd2889, 16'd16746, 16'd18470, 16'd57005, 16'd41078, 16'd55831}; // indx = 1872
    #10;
    addra = 32'd59936;
    dina = {96'd0, 16'd47074, 16'd64775, 16'd7833, 16'd25615, 16'd1523, 16'd28466, 16'd14835, 16'd61124, 16'd52181, 16'd54561}; // indx = 1873
    #10;
    addra = 32'd59968;
    dina = {96'd0, 16'd26893, 16'd60437, 16'd7707, 16'd56815, 16'd16819, 16'd35919, 16'd45867, 16'd44326, 16'd12888, 16'd24965}; // indx = 1874
    #10;
    addra = 32'd60000;
    dina = {96'd0, 16'd28570, 16'd35915, 16'd57850, 16'd62587, 16'd42947, 16'd42402, 16'd59825, 16'd5020, 16'd44050, 16'd24412}; // indx = 1875
    #10;
    addra = 32'd60032;
    dina = {96'd0, 16'd45959, 16'd1114, 16'd43279, 16'd32769, 16'd45527, 16'd26634, 16'd23927, 16'd28708, 16'd7631, 16'd11312}; // indx = 1876
    #10;
    addra = 32'd60064;
    dina = {96'd0, 16'd21917, 16'd24910, 16'd28456, 16'd57845, 16'd48262, 16'd62706, 16'd57091, 16'd14058, 16'd52754, 16'd20783}; // indx = 1877
    #10;
    addra = 32'd60096;
    dina = {96'd0, 16'd45859, 16'd39022, 16'd12162, 16'd39413, 16'd6333, 16'd49674, 16'd37475, 16'd59027, 16'd26804, 16'd31800}; // indx = 1878
    #10;
    addra = 32'd60128;
    dina = {96'd0, 16'd16154, 16'd56886, 16'd10962, 16'd7111, 16'd40902, 16'd6727, 16'd3409, 16'd28185, 16'd30485, 16'd12003}; // indx = 1879
    #10;
    addra = 32'd60160;
    dina = {96'd0, 16'd17394, 16'd45433, 16'd2233, 16'd47286, 16'd41655, 16'd1902, 16'd3305, 16'd58156, 16'd62518, 16'd5824}; // indx = 1880
    #10;
    addra = 32'd60192;
    dina = {96'd0, 16'd2188, 16'd382, 16'd64263, 16'd13263, 16'd36681, 16'd11922, 16'd28154, 16'd62313, 16'd9025, 16'd48798}; // indx = 1881
    #10;
    addra = 32'd60224;
    dina = {96'd0, 16'd46874, 16'd13132, 16'd33733, 16'd14748, 16'd29163, 16'd37765, 16'd31672, 16'd8391, 16'd38851, 16'd35163}; // indx = 1882
    #10;
    addra = 32'd60256;
    dina = {96'd0, 16'd24393, 16'd55111, 16'd59009, 16'd13433, 16'd3144, 16'd59401, 16'd62694, 16'd22151, 16'd53264, 16'd61307}; // indx = 1883
    #10;
    addra = 32'd60288;
    dina = {96'd0, 16'd49911, 16'd38788, 16'd12286, 16'd20375, 16'd5241, 16'd65016, 16'd16928, 16'd37354, 16'd36497, 16'd18613}; // indx = 1884
    #10;
    addra = 32'd60320;
    dina = {96'd0, 16'd18675, 16'd47397, 16'd9683, 16'd36037, 16'd2047, 16'd37807, 16'd46757, 16'd25374, 16'd50273, 16'd51950}; // indx = 1885
    #10;
    addra = 32'd60352;
    dina = {96'd0, 16'd15555, 16'd29449, 16'd48431, 16'd38894, 16'd11637, 16'd20983, 16'd16934, 16'd27961, 16'd34988, 16'd65257}; // indx = 1886
    #10;
    addra = 32'd60384;
    dina = {96'd0, 16'd11469, 16'd110, 16'd30918, 16'd9964, 16'd6860, 16'd44841, 16'd35397, 16'd14204, 16'd61613, 16'd10107}; // indx = 1887
    #10;
    addra = 32'd60416;
    dina = {96'd0, 16'd9343, 16'd51178, 16'd16580, 16'd25151, 16'd50650, 16'd27617, 16'd44942, 16'd11572, 16'd36069, 16'd16290}; // indx = 1888
    #10;
    addra = 32'd60448;
    dina = {96'd0, 16'd52618, 16'd38733, 16'd61543, 16'd50619, 16'd40088, 16'd6959, 16'd29925, 16'd63539, 16'd16588, 16'd33981}; // indx = 1889
    #10;
    addra = 32'd60480;
    dina = {96'd0, 16'd52438, 16'd29106, 16'd9046, 16'd52292, 16'd43117, 16'd63362, 16'd40826, 16'd52095, 16'd50281, 16'd21972}; // indx = 1890
    #10;
    addra = 32'd60512;
    dina = {96'd0, 16'd61357, 16'd16817, 16'd63154, 16'd18646, 16'd42638, 16'd64475, 16'd409, 16'd12929, 16'd56686, 16'd30107}; // indx = 1891
    #10;
    addra = 32'd60544;
    dina = {96'd0, 16'd2627, 16'd4379, 16'd23369, 16'd21478, 16'd7145, 16'd7651, 16'd15183, 16'd44513, 16'd29183, 16'd55318}; // indx = 1892
    #10;
    addra = 32'd60576;
    dina = {96'd0, 16'd52888, 16'd10156, 16'd12427, 16'd39871, 16'd22467, 16'd38756, 16'd13057, 16'd56096, 16'd45975, 16'd46536}; // indx = 1893
    #10;
    addra = 32'd60608;
    dina = {96'd0, 16'd11972, 16'd56958, 16'd16222, 16'd22550, 16'd14212, 16'd19239, 16'd11594, 16'd45627, 16'd16250, 16'd21161}; // indx = 1894
    #10;
    addra = 32'd60640;
    dina = {96'd0, 16'd40010, 16'd36531, 16'd61299, 16'd21251, 16'd60370, 16'd3867, 16'd1376, 16'd14183, 16'd13039, 16'd43273}; // indx = 1895
    #10;
    addra = 32'd60672;
    dina = {96'd0, 16'd59991, 16'd63851, 16'd2739, 16'd23599, 16'd31950, 16'd10989, 16'd30808, 16'd40318, 16'd21681, 16'd45276}; // indx = 1896
    #10;
    addra = 32'd60704;
    dina = {96'd0, 16'd43636, 16'd42184, 16'd2037, 16'd34428, 16'd20546, 16'd36203, 16'd42762, 16'd64590, 16'd54406, 16'd40747}; // indx = 1897
    #10;
    addra = 32'd60736;
    dina = {96'd0, 16'd18072, 16'd56303, 16'd9128, 16'd3371, 16'd26718, 16'd53544, 16'd5158, 16'd57233, 16'd61992, 16'd35829}; // indx = 1898
    #10;
    addra = 32'd60768;
    dina = {96'd0, 16'd29743, 16'd35589, 16'd56527, 16'd18784, 16'd49230, 16'd4976, 16'd16873, 16'd32640, 16'd26969, 16'd36334}; // indx = 1899
    #10;
    addra = 32'd60800;
    dina = {96'd0, 16'd46298, 16'd37124, 16'd21401, 16'd13280, 16'd50047, 16'd59838, 16'd29151, 16'd45597, 16'd4559, 16'd7332}; // indx = 1900
    #10;
    addra = 32'd60832;
    dina = {96'd0, 16'd9852, 16'd43890, 16'd35134, 16'd44105, 16'd4825, 16'd11290, 16'd44248, 16'd10043, 16'd12647, 16'd29517}; // indx = 1901
    #10;
    addra = 32'd60864;
    dina = {96'd0, 16'd22693, 16'd51661, 16'd19507, 16'd34967, 16'd34798, 16'd65311, 16'd12682, 16'd54613, 16'd22455, 16'd19862}; // indx = 1902
    #10;
    addra = 32'd60896;
    dina = {96'd0, 16'd56890, 16'd59903, 16'd25588, 16'd45822, 16'd36168, 16'd13701, 16'd13534, 16'd2779, 16'd3729, 16'd193}; // indx = 1903
    #10;
    addra = 32'd60928;
    dina = {96'd0, 16'd25348, 16'd28814, 16'd28420, 16'd28365, 16'd9361, 16'd2617, 16'd42313, 16'd61538, 16'd33186, 16'd50649}; // indx = 1904
    #10;
    addra = 32'd60960;
    dina = {96'd0, 16'd1800, 16'd47977, 16'd44085, 16'd12295, 16'd28813, 16'd49099, 16'd22045, 16'd14678, 16'd6287, 16'd36674}; // indx = 1905
    #10;
    addra = 32'd60992;
    dina = {96'd0, 16'd64558, 16'd35715, 16'd32426, 16'd19042, 16'd32389, 16'd11293, 16'd61425, 16'd58768, 16'd9536, 16'd41907}; // indx = 1906
    #10;
    addra = 32'd61024;
    dina = {96'd0, 16'd35303, 16'd58718, 16'd32255, 16'd27845, 16'd36165, 16'd18868, 16'd16659, 16'd9550, 16'd54132, 16'd49449}; // indx = 1907
    #10;
    addra = 32'd61056;
    dina = {96'd0, 16'd49604, 16'd16141, 16'd52310, 16'd19916, 16'd2542, 16'd30783, 16'd520, 16'd47075, 16'd64721, 16'd25615}; // indx = 1908
    #10;
    addra = 32'd61088;
    dina = {96'd0, 16'd55276, 16'd27039, 16'd25672, 16'd53087, 16'd55069, 16'd30396, 16'd13184, 16'd22933, 16'd16694, 16'd5157}; // indx = 1909
    #10;
    addra = 32'd61120;
    dina = {96'd0, 16'd13950, 16'd11543, 16'd20794, 16'd13561, 16'd35267, 16'd32991, 16'd20637, 16'd59759, 16'd46733, 16'd56710}; // indx = 1910
    #10;
    addra = 32'd61152;
    dina = {96'd0, 16'd21374, 16'd19261, 16'd31947, 16'd40156, 16'd28837, 16'd23716, 16'd42499, 16'd22615, 16'd48441, 16'd23097}; // indx = 1911
    #10;
    addra = 32'd61184;
    dina = {96'd0, 16'd55956, 16'd26426, 16'd17745, 16'd24039, 16'd59569, 16'd53013, 16'd35551, 16'd40758, 16'd30242, 16'd55794}; // indx = 1912
    #10;
    addra = 32'd61216;
    dina = {96'd0, 16'd51885, 16'd2375, 16'd29827, 16'd64400, 16'd61420, 16'd56751, 16'd36388, 16'd12429, 16'd38587, 16'd54075}; // indx = 1913
    #10;
    addra = 32'd61248;
    dina = {96'd0, 16'd7136, 16'd32733, 16'd48122, 16'd46350, 16'd34159, 16'd5292, 16'd47904, 16'd15643, 16'd8586, 16'd29442}; // indx = 1914
    #10;
    addra = 32'd61280;
    dina = {96'd0, 16'd16143, 16'd30061, 16'd31814, 16'd21301, 16'd8562, 16'd62337, 16'd125, 16'd52883, 16'd6479, 16'd40056}; // indx = 1915
    #10;
    addra = 32'd61312;
    dina = {96'd0, 16'd44796, 16'd1024, 16'd32845, 16'd34960, 16'd5579, 16'd47410, 16'd61678, 16'd26186, 16'd21114, 16'd2325}; // indx = 1916
    #10;
    addra = 32'd61344;
    dina = {96'd0, 16'd30398, 16'd29184, 16'd24556, 16'd6328, 16'd57278, 16'd44515, 16'd53875, 16'd26941, 16'd3506, 16'd45561}; // indx = 1917
    #10;
    addra = 32'd61376;
    dina = {96'd0, 16'd52301, 16'd20571, 16'd2914, 16'd64149, 16'd11549, 16'd27410, 16'd17416, 16'd24298, 16'd58987, 16'd54586}; // indx = 1918
    #10;
    addra = 32'd61408;
    dina = {96'd0, 16'd61137, 16'd53172, 16'd9339, 16'd12345, 16'd12772, 16'd30743, 16'd41443, 16'd22361, 16'd65433, 16'd42177}; // indx = 1919
    #10;
    addra = 32'd61440;
    dina = {96'd0, 16'd40052, 16'd21235, 16'd23394, 16'd49397, 16'd9402, 16'd56856, 16'd61432, 16'd13116, 16'd52558, 16'd19509}; // indx = 1920
    #10;
    addra = 32'd61472;
    dina = {96'd0, 16'd40282, 16'd3856, 16'd4355, 16'd27913, 16'd10781, 16'd2408, 16'd17599, 16'd12036, 16'd56353, 16'd15133}; // indx = 1921
    #10;
    addra = 32'd61504;
    dina = {96'd0, 16'd8979, 16'd235, 16'd22071, 16'd30388, 16'd22474, 16'd42577, 16'd26200, 16'd27603, 16'd10953, 16'd25335}; // indx = 1922
    #10;
    addra = 32'd61536;
    dina = {96'd0, 16'd33982, 16'd42297, 16'd677, 16'd54293, 16'd28647, 16'd15509, 16'd28626, 16'd63156, 16'd14980, 16'd9032}; // indx = 1923
    #10;
    addra = 32'd61568;
    dina = {96'd0, 16'd63705, 16'd50250, 16'd25072, 16'd63282, 16'd3043, 16'd15865, 16'd18584, 16'd48364, 16'd24370, 16'd34056}; // indx = 1924
    #10;
    addra = 32'd61600;
    dina = {96'd0, 16'd16327, 16'd3437, 16'd58271, 16'd49079, 16'd4375, 16'd25905, 16'd8739, 16'd31516, 16'd58599, 16'd26878}; // indx = 1925
    #10;
    addra = 32'd61632;
    dina = {96'd0, 16'd11395, 16'd42566, 16'd25861, 16'd34187, 16'd33638, 16'd58808, 16'd8727, 16'd12570, 16'd25895, 16'd22383}; // indx = 1926
    #10;
    addra = 32'd61664;
    dina = {96'd0, 16'd36914, 16'd43197, 16'd26937, 16'd42679, 16'd61754, 16'd39940, 16'd63856, 16'd38072, 16'd55418, 16'd65488}; // indx = 1927
    #10;
    addra = 32'd61696;
    dina = {96'd0, 16'd43344, 16'd46018, 16'd17237, 16'd18041, 16'd26433, 16'd19738, 16'd15528, 16'd33201, 16'd62859, 16'd12455}; // indx = 1928
    #10;
    addra = 32'd61728;
    dina = {96'd0, 16'd34792, 16'd15254, 16'd7833, 16'd51683, 16'd24748, 16'd21275, 16'd3891, 16'd62957, 16'd49948, 16'd40704}; // indx = 1929
    #10;
    addra = 32'd61760;
    dina = {96'd0, 16'd34051, 16'd28637, 16'd23495, 16'd27764, 16'd57092, 16'd44090, 16'd1274, 16'd780, 16'd27823, 16'd25870}; // indx = 1930
    #10;
    addra = 32'd61792;
    dina = {96'd0, 16'd22682, 16'd25108, 16'd45764, 16'd53809, 16'd30059, 16'd64436, 16'd25730, 16'd1811, 16'd43740, 16'd9910}; // indx = 1931
    #10;
    addra = 32'd61824;
    dina = {96'd0, 16'd38439, 16'd22168, 16'd31831, 16'd62181, 16'd43945, 16'd53954, 16'd36119, 16'd40372, 16'd53654, 16'd17372}; // indx = 1932
    #10;
    addra = 32'd61856;
    dina = {96'd0, 16'd58756, 16'd25273, 16'd18959, 16'd32456, 16'd47244, 16'd20552, 16'd52369, 16'd26103, 16'd41273, 16'd19713}; // indx = 1933
    #10;
    addra = 32'd61888;
    dina = {96'd0, 16'd23617, 16'd24450, 16'd37669, 16'd33773, 16'd34543, 16'd21522, 16'd58654, 16'd18319, 16'd51962, 16'd17447}; // indx = 1934
    #10;
    addra = 32'd61920;
    dina = {96'd0, 16'd44665, 16'd10905, 16'd56671, 16'd20282, 16'd43909, 16'd7800, 16'd57950, 16'd17805, 16'd30782, 16'd29663}; // indx = 1935
    #10;
    addra = 32'd61952;
    dina = {96'd0, 16'd53012, 16'd26345, 16'd16909, 16'd28091, 16'd49048, 16'd16609, 16'd46914, 16'd8550, 16'd34052, 16'd48261}; // indx = 1936
    #10;
    addra = 32'd61984;
    dina = {96'd0, 16'd30063, 16'd18532, 16'd3871, 16'd46243, 16'd57259, 16'd10893, 16'd4187, 16'd3160, 16'd7135, 16'd23930}; // indx = 1937
    #10;
    addra = 32'd62016;
    dina = {96'd0, 16'd1005, 16'd20313, 16'd43291, 16'd46925, 16'd21096, 16'd43792, 16'd15612, 16'd55976, 16'd826, 16'd26476}; // indx = 1938
    #10;
    addra = 32'd62048;
    dina = {96'd0, 16'd52153, 16'd42783, 16'd61828, 16'd17323, 16'd27628, 16'd16919, 16'd21096, 16'd53368, 16'd36080, 16'd38703}; // indx = 1939
    #10;
    addra = 32'd62080;
    dina = {96'd0, 16'd63535, 16'd25004, 16'd44019, 16'd53525, 16'd33720, 16'd53004, 16'd22231, 16'd16269, 16'd14071, 16'd63718}; // indx = 1940
    #10;
    addra = 32'd62112;
    dina = {96'd0, 16'd58038, 16'd36290, 16'd6642, 16'd27950, 16'd10464, 16'd25812, 16'd45596, 16'd37082, 16'd53102, 16'd62548}; // indx = 1941
    #10;
    addra = 32'd62144;
    dina = {96'd0, 16'd30599, 16'd18597, 16'd12954, 16'd448, 16'd12665, 16'd60, 16'd14195, 16'd43162, 16'd35325, 16'd30835}; // indx = 1942
    #10;
    addra = 32'd62176;
    dina = {96'd0, 16'd43426, 16'd134, 16'd37912, 16'd58294, 16'd10008, 16'd4770, 16'd1846, 16'd42109, 16'd61139, 16'd55957}; // indx = 1943
    #10;
    addra = 32'd62208;
    dina = {96'd0, 16'd9572, 16'd60534, 16'd52251, 16'd14860, 16'd64158, 16'd29381, 16'd41454, 16'd40221, 16'd12695, 16'd46943}; // indx = 1944
    #10;
    addra = 32'd62240;
    dina = {96'd0, 16'd51061, 16'd54798, 16'd17958, 16'd30501, 16'd35277, 16'd38018, 16'd35524, 16'd18836, 16'd47573, 16'd5292}; // indx = 1945
    #10;
    addra = 32'd62272;
    dina = {96'd0, 16'd33698, 16'd22378, 16'd3016, 16'd19028, 16'd46859, 16'd21552, 16'd33086, 16'd26091, 16'd43436, 16'd62777}; // indx = 1946
    #10;
    addra = 32'd62304;
    dina = {96'd0, 16'd46521, 16'd1767, 16'd15202, 16'd8095, 16'd7452, 16'd37556, 16'd25412, 16'd58008, 16'd42366, 16'd78}; // indx = 1947
    #10;
    addra = 32'd62336;
    dina = {96'd0, 16'd31540, 16'd36288, 16'd25843, 16'd16274, 16'd59963, 16'd30556, 16'd61127, 16'd6109, 16'd32581, 16'd23994}; // indx = 1948
    #10;
    addra = 32'd62368;
    dina = {96'd0, 16'd29010, 16'd44487, 16'd12677, 16'd27423, 16'd45979, 16'd60631, 16'd51136, 16'd7639, 16'd35042, 16'd6469}; // indx = 1949
    #10;
    addra = 32'd62400;
    dina = {96'd0, 16'd542, 16'd39142, 16'd10516, 16'd43794, 16'd14312, 16'd52977, 16'd49164, 16'd8398, 16'd35668, 16'd17031}; // indx = 1950
    #10;
    addra = 32'd62432;
    dina = {96'd0, 16'd28910, 16'd56162, 16'd9377, 16'd16677, 16'd36413, 16'd26693, 16'd25912, 16'd63501, 16'd57026, 16'd35419}; // indx = 1951
    #10;
    addra = 32'd62464;
    dina = {96'd0, 16'd7972, 16'd13825, 16'd29193, 16'd44817, 16'd56947, 16'd45756, 16'd2298, 16'd21749, 16'd55464, 16'd60046}; // indx = 1952
    #10;
    addra = 32'd62496;
    dina = {96'd0, 16'd20832, 16'd27860, 16'd6887, 16'd33255, 16'd59766, 16'd28989, 16'd51896, 16'd12427, 16'd12603, 16'd20368}; // indx = 1953
    #10;
    addra = 32'd62528;
    dina = {96'd0, 16'd55035, 16'd15085, 16'd63472, 16'd209, 16'd29758, 16'd34169, 16'd53910, 16'd14608, 16'd19496, 16'd41063}; // indx = 1954
    #10;
    addra = 32'd62560;
    dina = {96'd0, 16'd38727, 16'd55418, 16'd30138, 16'd27336, 16'd35260, 16'd6422, 16'd63912, 16'd56310, 16'd30397, 16'd1940}; // indx = 1955
    #10;
    addra = 32'd62592;
    dina = {96'd0, 16'd60830, 16'd41013, 16'd1498, 16'd46261, 16'd13830, 16'd2591, 16'd10178, 16'd46769, 16'd64013, 16'd60557}; // indx = 1956
    #10;
    addra = 32'd62624;
    dina = {96'd0, 16'd9750, 16'd24266, 16'd21596, 16'd7151, 16'd56821, 16'd50850, 16'd4852, 16'd2349, 16'd39994, 16'd42018}; // indx = 1957
    #10;
    addra = 32'd62656;
    dina = {96'd0, 16'd16801, 16'd1666, 16'd27791, 16'd60862, 16'd51998, 16'd50753, 16'd55457, 16'd11898, 16'd21669, 16'd46765}; // indx = 1958
    #10;
    addra = 32'd62688;
    dina = {96'd0, 16'd26302, 16'd40966, 16'd29569, 16'd529, 16'd43986, 16'd44046, 16'd1691, 16'd25587, 16'd7325, 16'd3172}; // indx = 1959
    #10;
    addra = 32'd62720;
    dina = {96'd0, 16'd18791, 16'd1162, 16'd64797, 16'd13171, 16'd28193, 16'd51879, 16'd8770, 16'd53955, 16'd38559, 16'd56080}; // indx = 1960
    #10;
    addra = 32'd62752;
    dina = {96'd0, 16'd34501, 16'd31111, 16'd2987, 16'd14560, 16'd46268, 16'd34998, 16'd37740, 16'd36258, 16'd4651, 16'd15171}; // indx = 1961
    #10;
    addra = 32'd62784;
    dina = {96'd0, 16'd55115, 16'd49886, 16'd43449, 16'd20918, 16'd1998, 16'd54897, 16'd60691, 16'd49885, 16'd53132, 16'd17186}; // indx = 1962
    #10;
    addra = 32'd62816;
    dina = {96'd0, 16'd759, 16'd64844, 16'd3866, 16'd47314, 16'd45728, 16'd3541, 16'd35105, 16'd10789, 16'd22162, 16'd56405}; // indx = 1963
    #10;
    addra = 32'd62848;
    dina = {96'd0, 16'd34322, 16'd61927, 16'd1001, 16'd20193, 16'd49480, 16'd12480, 16'd17245, 16'd16811, 16'd15827, 16'd35946}; // indx = 1964
    #10;
    addra = 32'd62880;
    dina = {96'd0, 16'd23556, 16'd6465, 16'd4997, 16'd16289, 16'd50057, 16'd32698, 16'd14437, 16'd48444, 16'd9243, 16'd33196}; // indx = 1965
    #10;
    addra = 32'd62912;
    dina = {96'd0, 16'd46497, 16'd26902, 16'd51179, 16'd10974, 16'd46233, 16'd6963, 16'd21556, 16'd62304, 16'd64791, 16'd8078}; // indx = 1966
    #10;
    addra = 32'd62944;
    dina = {96'd0, 16'd35666, 16'd42144, 16'd50452, 16'd59306, 16'd41790, 16'd13217, 16'd45457, 16'd22760, 16'd12919, 16'd40762}; // indx = 1967
    #10;
    addra = 32'd62976;
    dina = {96'd0, 16'd37152, 16'd53942, 16'd50857, 16'd63354, 16'd55400, 16'd192, 16'd39233, 16'd60799, 16'd5252, 16'd17174}; // indx = 1968
    #10;
    addra = 32'd63008;
    dina = {96'd0, 16'd30063, 16'd51580, 16'd58972, 16'd30893, 16'd5516, 16'd2810, 16'd34670, 16'd65174, 16'd62394, 16'd35874}; // indx = 1969
    #10;
    addra = 32'd63040;
    dina = {96'd0, 16'd10527, 16'd62467, 16'd60489, 16'd64224, 16'd60117, 16'd14628, 16'd22000, 16'd8444, 16'd43904, 16'd6663}; // indx = 1970
    #10;
    addra = 32'd63072;
    dina = {96'd0, 16'd16673, 16'd28519, 16'd43315, 16'd15934, 16'd20344, 16'd54256, 16'd23673, 16'd56608, 16'd61106, 16'd19630}; // indx = 1971
    #10;
    addra = 32'd63104;
    dina = {96'd0, 16'd14604, 16'd56623, 16'd18424, 16'd1146, 16'd50334, 16'd10793, 16'd48674, 16'd53269, 16'd58740, 16'd45828}; // indx = 1972
    #10;
    addra = 32'd63136;
    dina = {96'd0, 16'd15860, 16'd56263, 16'd8644, 16'd28823, 16'd13189, 16'd43029, 16'd46455, 16'd42124, 16'd27065, 16'd10401}; // indx = 1973
    #10;
    addra = 32'd63168;
    dina = {96'd0, 16'd28565, 16'd39840, 16'd2748, 16'd2823, 16'd63209, 16'd24675, 16'd48805, 16'd9276, 16'd49965, 16'd54098}; // indx = 1974
    #10;
    addra = 32'd63200;
    dina = {96'd0, 16'd16386, 16'd50122, 16'd29222, 16'd24351, 16'd34017, 16'd50845, 16'd24629, 16'd867, 16'd44542, 16'd37318}; // indx = 1975
    #10;
    addra = 32'd63232;
    dina = {96'd0, 16'd17745, 16'd25931, 16'd52086, 16'd4527, 16'd16041, 16'd19710, 16'd44663, 16'd13948, 16'd5072, 16'd42025}; // indx = 1976
    #10;
    addra = 32'd63264;
    dina = {96'd0, 16'd1451, 16'd56417, 16'd9770, 16'd10647, 16'd24743, 16'd19477, 16'd46409, 16'd64353, 16'd42167, 16'd26803}; // indx = 1977
    #10;
    addra = 32'd63296;
    dina = {96'd0, 16'd7840, 16'd3146, 16'd56881, 16'd52518, 16'd26188, 16'd23126, 16'd33259, 16'd55455, 16'd16630, 16'd2754}; // indx = 1978
    #10;
    addra = 32'd63328;
    dina = {96'd0, 16'd30889, 16'd18069, 16'd8369, 16'd6881, 16'd9168, 16'd14535, 16'd31720, 16'd1788, 16'd54780, 16'd30808}; // indx = 1979
    #10;
    addra = 32'd63360;
    dina = {96'd0, 16'd43430, 16'd11996, 16'd9127, 16'd994, 16'd61594, 16'd14692, 16'd14848, 16'd20882, 16'd15271, 16'd12569}; // indx = 1980
    #10;
    addra = 32'd63392;
    dina = {96'd0, 16'd39485, 16'd6005, 16'd4387, 16'd64997, 16'd31836, 16'd56895, 16'd37676, 16'd15229, 16'd11881, 16'd54623}; // indx = 1981
    #10;
    addra = 32'd63424;
    dina = {96'd0, 16'd42410, 16'd24921, 16'd51211, 16'd46895, 16'd64684, 16'd46992, 16'd61062, 16'd33064, 16'd57940, 16'd8053}; // indx = 1982
    #10;
    addra = 32'd63456;
    dina = {96'd0, 16'd16576, 16'd60122, 16'd11082, 16'd5205, 16'd5514, 16'd12915, 16'd58698, 16'd62596, 16'd18525, 16'd64009}; // indx = 1983
    #10;
    addra = 32'd63488;
    dina = {96'd0, 16'd11078, 16'd54949, 16'd64684, 16'd10207, 16'd36661, 16'd51821, 16'd31397, 16'd44578, 16'd38753, 16'd669}; // indx = 1984
    #10;
    addra = 32'd63520;
    dina = {96'd0, 16'd48038, 16'd19661, 16'd22114, 16'd54767, 16'd64327, 16'd14949, 16'd29784, 16'd34011, 16'd45203, 16'd47766}; // indx = 1985
    #10;
    addra = 32'd63552;
    dina = {96'd0, 16'd12148, 16'd43142, 16'd6095, 16'd35008, 16'd31064, 16'd10076, 16'd15825, 16'd45452, 16'd38258, 16'd8971}; // indx = 1986
    #10;
    addra = 32'd63584;
    dina = {96'd0, 16'd22108, 16'd57330, 16'd13783, 16'd4829, 16'd43601, 16'd5518, 16'd47373, 16'd19206, 16'd6434, 16'd5075}; // indx = 1987
    #10;
    addra = 32'd63616;
    dina = {96'd0, 16'd20177, 16'd49451, 16'd21186, 16'd21533, 16'd52391, 16'd51754, 16'd5231, 16'd19426, 16'd30589, 16'd833}; // indx = 1988
    #10;
    addra = 32'd63648;
    dina = {96'd0, 16'd50585, 16'd384, 16'd14436, 16'd6255, 16'd11796, 16'd60607, 16'd47922, 16'd60407, 16'd7564, 16'd5602}; // indx = 1989
    #10;
    addra = 32'd63680;
    dina = {96'd0, 16'd52093, 16'd55954, 16'd6994, 16'd32450, 16'd310, 16'd3434, 16'd6671, 16'd34686, 16'd39635, 16'd17678}; // indx = 1990
    #10;
    addra = 32'd63712;
    dina = {96'd0, 16'd2250, 16'd52666, 16'd28893, 16'd20913, 16'd8602, 16'd18241, 16'd43773, 16'd57668, 16'd51472, 16'd19488}; // indx = 1991
    #10;
    addra = 32'd63744;
    dina = {96'd0, 16'd29185, 16'd30788, 16'd41977, 16'd41890, 16'd7082, 16'd30629, 16'd7321, 16'd42574, 16'd7052, 16'd30940}; // indx = 1992
    #10;
    addra = 32'd63776;
    dina = {96'd0, 16'd49345, 16'd8617, 16'd29587, 16'd39071, 16'd56810, 16'd57349, 16'd54105, 16'd48821, 16'd22627, 16'd39948}; // indx = 1993
    #10;
    addra = 32'd63808;
    dina = {96'd0, 16'd11847, 16'd14231, 16'd49599, 16'd38473, 16'd10381, 16'd24029, 16'd1315, 16'd3778, 16'd29480, 16'd28300}; // indx = 1994
    #10;
    addra = 32'd63840;
    dina = {96'd0, 16'd54985, 16'd25991, 16'd10563, 16'd32090, 16'd29409, 16'd19397, 16'd9661, 16'd58988, 16'd48835, 16'd21592}; // indx = 1995
    #10;
    addra = 32'd63872;
    dina = {96'd0, 16'd14034, 16'd46137, 16'd9758, 16'd52835, 16'd41805, 16'd42576, 16'd9232, 16'd59605, 16'd18791, 16'd26423}; // indx = 1996
    #10;
    addra = 32'd63904;
    dina = {96'd0, 16'd24272, 16'd12912, 16'd19047, 16'd49669, 16'd24276, 16'd13076, 16'd43084, 16'd31152, 16'd4401, 16'd32075}; // indx = 1997
    #10;
    addra = 32'd63936;
    dina = {96'd0, 16'd10047, 16'd62858, 16'd61855, 16'd28125, 16'd21628, 16'd27854, 16'd15511, 16'd10989, 16'd22261, 16'd44448}; // indx = 1998
    #10;
    addra = 32'd63968;
    dina = {96'd0, 16'd10122, 16'd3142, 16'd46910, 16'd24278, 16'd60369, 16'd52181, 16'd1652, 16'd7597, 16'd12725, 16'd33098}; // indx = 1999
    #10;
    addra = 32'd64000;
    dina = {96'd0, 16'd2512, 16'd9886, 16'd16073, 16'd23917, 16'd31829, 16'd444, 16'd14432, 16'd46406, 16'd16966, 16'd49961}; // indx = 2000
    #10;
    addra = 32'd64032;
    dina = {96'd0, 16'd9555, 16'd8669, 16'd60541, 16'd61506, 16'd49521, 16'd61214, 16'd4571, 16'd31721, 16'd48492, 16'd18800}; // indx = 2001
    #10;
    addra = 32'd64064;
    dina = {96'd0, 16'd7665, 16'd26243, 16'd14298, 16'd53396, 16'd32467, 16'd12605, 16'd49437, 16'd3803, 16'd7965, 16'd13762}; // indx = 2002
    #10;
    addra = 32'd64096;
    dina = {96'd0, 16'd21418, 16'd42657, 16'd45467, 16'd14013, 16'd16620, 16'd53426, 16'd59284, 16'd25324, 16'd12621, 16'd33880}; // indx = 2003
    #10;
    addra = 32'd64128;
    dina = {96'd0, 16'd19424, 16'd33858, 16'd23953, 16'd44963, 16'd7235, 16'd57964, 16'd132, 16'd43228, 16'd1012, 16'd28591}; // indx = 2004
    #10;
    addra = 32'd64160;
    dina = {96'd0, 16'd6867, 16'd14266, 16'd56577, 16'd9032, 16'd6151, 16'd36867, 16'd34099, 16'd6755, 16'd10847, 16'd20431}; // indx = 2005
    #10;
    addra = 32'd64192;
    dina = {96'd0, 16'd57361, 16'd28455, 16'd25782, 16'd34942, 16'd62803, 16'd55345, 16'd33118, 16'd58247, 16'd5156, 16'd57449}; // indx = 2006
    #10;
    addra = 32'd64224;
    dina = {96'd0, 16'd29921, 16'd49940, 16'd53537, 16'd19033, 16'd50679, 16'd60639, 16'd11882, 16'd18820, 16'd55229, 16'd9915}; // indx = 2007
    #10;
    addra = 32'd64256;
    dina = {96'd0, 16'd48268, 16'd59265, 16'd24078, 16'd51739, 16'd5450, 16'd6949, 16'd49364, 16'd54796, 16'd55442, 16'd14204}; // indx = 2008
    #10;
    addra = 32'd64288;
    dina = {96'd0, 16'd19754, 16'd28280, 16'd63282, 16'd52365, 16'd37430, 16'd58996, 16'd10737, 16'd59167, 16'd8417, 16'd57162}; // indx = 2009
    #10;
    addra = 32'd64320;
    dina = {96'd0, 16'd55346, 16'd6989, 16'd26944, 16'd28358, 16'd56733, 16'd9245, 16'd6091, 16'd14851, 16'd15832, 16'd10550}; // indx = 2010
    #10;
    addra = 32'd64352;
    dina = {96'd0, 16'd35831, 16'd15104, 16'd48933, 16'd17459, 16'd29919, 16'd32367, 16'd32907, 16'd12236, 16'd31697, 16'd29616}; // indx = 2011
    #10;
    addra = 32'd64384;
    dina = {96'd0, 16'd25452, 16'd34154, 16'd38573, 16'd27035, 16'd26780, 16'd38756, 16'd8308, 16'd17413, 16'd49087, 16'd38356}; // indx = 2012
    #10;
    addra = 32'd64416;
    dina = {96'd0, 16'd63220, 16'd51714, 16'd11557, 16'd45459, 16'd665, 16'd4928, 16'd19118, 16'd14535, 16'd52846, 16'd12715}; // indx = 2013
    #10;
    addra = 32'd64448;
    dina = {96'd0, 16'd18403, 16'd22715, 16'd16788, 16'd37086, 16'd55796, 16'd8128, 16'd21710, 16'd27102, 16'd7605, 16'd33294}; // indx = 2014
    #10;
    addra = 32'd64480;
    dina = {96'd0, 16'd1611, 16'd24470, 16'd26106, 16'd19322, 16'd35376, 16'd54166, 16'd19064, 16'd35699, 16'd46021, 16'd54246}; // indx = 2015
    #10;
    addra = 32'd64512;
    dina = {96'd0, 16'd49901, 16'd7280, 16'd8954, 16'd18849, 16'd34222, 16'd313, 16'd4795, 16'd61640, 16'd58832, 16'd9818}; // indx = 2016
    #10;
    addra = 32'd64544;
    dina = {96'd0, 16'd19862, 16'd6912, 16'd8243, 16'd55991, 16'd8693, 16'd62905, 16'd58633, 16'd37114, 16'd37537, 16'd54838}; // indx = 2017
    #10;
    addra = 32'd64576;
    dina = {96'd0, 16'd51859, 16'd37857, 16'd58328, 16'd48737, 16'd1311, 16'd26017, 16'd15220, 16'd5726, 16'd30740, 16'd5679}; // indx = 2018
    #10;
    addra = 32'd64608;
    dina = {96'd0, 16'd41962, 16'd15141, 16'd33183, 16'd6012, 16'd21144, 16'd32736, 16'd32266, 16'd31672, 16'd24035, 16'd23508}; // indx = 2019
    #10;
    addra = 32'd64640;
    dina = {96'd0, 16'd43664, 16'd44475, 16'd34509, 16'd22813, 16'd5145, 16'd63311, 16'd37866, 16'd37457, 16'd25085, 16'd736}; // indx = 2020
    #10;
    addra = 32'd64672;
    dina = {96'd0, 16'd42488, 16'd7903, 16'd18856, 16'd52403, 16'd34840, 16'd40687, 16'd46428, 16'd24371, 16'd9123, 16'd22887}; // indx = 2021
    #10;
    addra = 32'd64704;
    dina = {96'd0, 16'd51210, 16'd1316, 16'd9414, 16'd50731, 16'd40299, 16'd39698, 16'd11534, 16'd33372, 16'd16700, 16'd39305}; // indx = 2022
    #10;
    addra = 32'd64736;
    dina = {96'd0, 16'd17113, 16'd37924, 16'd58822, 16'd7461, 16'd56742, 16'd57364, 16'd55048, 16'd57545, 16'd34545, 16'd33207}; // indx = 2023
    #10;
    addra = 32'd64768;
    dina = {96'd0, 16'd52730, 16'd6518, 16'd38667, 16'd44177, 16'd64573, 16'd34079, 16'd19988, 16'd7309, 16'd17139, 16'd46196}; // indx = 2024
    #10;
    addra = 32'd64800;
    dina = {96'd0, 16'd52333, 16'd13298, 16'd6123, 16'd16672, 16'd6183, 16'd22147, 16'd50459, 16'd20292, 16'd62877, 16'd58659}; // indx = 2025
    #10;
    addra = 32'd64832;
    dina = {96'd0, 16'd56766, 16'd22788, 16'd55742, 16'd16029, 16'd33351, 16'd927, 16'd18960, 16'd17802, 16'd60707, 16'd4722}; // indx = 2026
    #10;
    addra = 32'd64864;
    dina = {96'd0, 16'd24359, 16'd19845, 16'd32331, 16'd45565, 16'd61188, 16'd34681, 16'd7083, 16'd46247, 16'd63542, 16'd48026}; // indx = 2027
    #10;
    addra = 32'd64896;
    dina = {96'd0, 16'd33314, 16'd24673, 16'd40463, 16'd64733, 16'd57717, 16'd33649, 16'd55479, 16'd35664, 16'd49453, 16'd45074}; // indx = 2028
    #10;
    addra = 32'd64928;
    dina = {96'd0, 16'd2861, 16'd46660, 16'd57765, 16'd28054, 16'd11076, 16'd38628, 16'd61677, 16'd34095, 16'd34127, 16'd14393}; // indx = 2029
    #10;
    addra = 32'd64960;
    dina = {96'd0, 16'd31203, 16'd8555, 16'd2954, 16'd21425, 16'd56968, 16'd56408, 16'd61263, 16'd18420, 16'd39367, 16'd34844}; // indx = 2030
    #10;
    addra = 32'd64992;
    dina = {96'd0, 16'd51961, 16'd12057, 16'd32347, 16'd57919, 16'd46377, 16'd14913, 16'd27111, 16'd10119, 16'd7190, 16'd60852}; // indx = 2031
    #10;
    addra = 32'd65024;
    dina = {96'd0, 16'd19177, 16'd34399, 16'd54822, 16'd25837, 16'd28487, 16'd4279, 16'd60623, 16'd53067, 16'd1860, 16'd57246}; // indx = 2032
    #10;
    addra = 32'd65056;
    dina = {96'd0, 16'd49991, 16'd18501, 16'd49458, 16'd3340, 16'd36357, 16'd20554, 16'd1915, 16'd31605, 16'd53468, 16'd15084}; // indx = 2033
    #10;
    addra = 32'd65088;
    dina = {96'd0, 16'd20575, 16'd15242, 16'd55523, 16'd43352, 16'd3113, 16'd5709, 16'd21137, 16'd53093, 16'd14418, 16'd30345}; // indx = 2034
    #10;
    addra = 32'd65120;
    dina = {96'd0, 16'd51741, 16'd58367, 16'd5262, 16'd23934, 16'd20366, 16'd57728, 16'd30424, 16'd62857, 16'd55863, 16'd21597}; // indx = 2035
    #10;
    addra = 32'd65152;
    dina = {96'd0, 16'd25976, 16'd9438, 16'd37441, 16'd15370, 16'd36902, 16'd28344, 16'd13546, 16'd3012, 16'd52243, 16'd49741}; // indx = 2036
    #10;
    addra = 32'd65184;
    dina = {96'd0, 16'd56797, 16'd4756, 16'd18628, 16'd54655, 16'd25991, 16'd50022, 16'd11175, 16'd36711, 16'd7688, 16'd17797}; // indx = 2037
    #10;
    addra = 32'd65216;
    dina = {96'd0, 16'd9170, 16'd50254, 16'd36560, 16'd25687, 16'd17324, 16'd54053, 16'd44177, 16'd58182, 16'd40222, 16'd55453}; // indx = 2038
    #10;
    addra = 32'd65248;
    dina = {96'd0, 16'd54436, 16'd49965, 16'd14144, 16'd8624, 16'd36431, 16'd22697, 16'd53514, 16'd63757, 16'd41986, 16'd29895}; // indx = 2039
    #10;
    addra = 32'd65280;
    dina = {96'd0, 16'd15044, 16'd32028, 16'd31063, 16'd32568, 16'd60529, 16'd25349, 16'd45119, 16'd47130, 16'd10162, 16'd29703}; // indx = 2040
    #10;
    addra = 32'd65312;
    dina = {96'd0, 16'd4582, 16'd18106, 16'd26716, 16'd17882, 16'd35975, 16'd56067, 16'd1513, 16'd11962, 16'd60218, 16'd16641}; // indx = 2041
    #10;
    addra = 32'd65344;
    dina = {96'd0, 16'd40319, 16'd3844, 16'd59478, 16'd11623, 16'd17215, 16'd37675, 16'd39489, 16'd27405, 16'd25655, 16'd31634}; // indx = 2042
    #10;
    addra = 32'd65376;
    dina = {96'd0, 16'd40935, 16'd62411, 16'd57044, 16'd44896, 16'd54079, 16'd4200, 16'd38304, 16'd27032, 16'd35760, 16'd64959}; // indx = 2043
    #10;
    addra = 32'd65408;
    dina = {96'd0, 16'd22573, 16'd7358, 16'd45685, 16'd548, 16'd32383, 16'd4558, 16'd34302, 16'd56231, 16'd50547, 16'd9102}; // indx = 2044
    #10;
    addra = 32'd65440;
    dina = {96'd0, 16'd2991, 16'd20141, 16'd55721, 16'd46741, 16'd22774, 16'd48533, 16'd1504, 16'd19230, 16'd44342, 16'd40502}; // indx = 2045
    #10;
    addra = 32'd65472;
    dina = {96'd0, 16'd65075, 16'd9079, 16'd39476, 16'd1710, 16'd44532, 16'd21562, 16'd53954, 16'd40583, 16'd3933, 16'd29945}; // indx = 2046
    #10;
    addra = 32'd65504;
    dina = {96'd0, 16'd34710, 16'd54016, 16'd42333, 16'd21534, 16'd13694, 16'd28132, 16'd28902, 16'd28007, 16'd59534, 16'd11316}; // indx = 2047
    #10;
    addra = 32'd65536;
    dina = {96'd0, 16'd50773, 16'd22207, 16'd16131, 16'd16827, 16'd56173, 16'd13549, 16'd59759, 16'd32089, 16'd1594, 16'd47435}; // indx = 2048
    #10;
    addra = 32'd65568;
    dina = {96'd0, 16'd56833, 16'd49040, 16'd14738, 16'd40451, 16'd41219, 16'd47152, 16'd10913, 16'd63326, 16'd3037, 16'd14003}; // indx = 2049
    #10;
    addra = 32'd65600;
    dina = {96'd0, 16'd32466, 16'd6707, 16'd56563, 16'd49065, 16'd29531, 16'd57301, 16'd18057, 16'd48183, 16'd54679, 16'd31881}; // indx = 2050
    #10;
    addra = 32'd65632;
    dina = {96'd0, 16'd61595, 16'd7324, 16'd57943, 16'd25721, 16'd54143, 16'd48571, 16'd36825, 16'd8735, 16'd46667, 16'd61230}; // indx = 2051
    #10;
    addra = 32'd65664;
    dina = {96'd0, 16'd21283, 16'd7874, 16'd43574, 16'd36209, 16'd12775, 16'd54396, 16'd32475, 16'd53670, 16'd25606, 16'd14751}; // indx = 2052
    #10;
    addra = 32'd65696;
    dina = {96'd0, 16'd60251, 16'd29712, 16'd13415, 16'd12668, 16'd13511, 16'd7231, 16'd20239, 16'd61060, 16'd18952, 16'd60647}; // indx = 2053
    #10;
    addra = 32'd65728;
    dina = {96'd0, 16'd31659, 16'd56585, 16'd31611, 16'd27995, 16'd7991, 16'd20220, 16'd19551, 16'd52440, 16'd29306, 16'd59145}; // indx = 2054
    #10;
    addra = 32'd65760;
    dina = {96'd0, 16'd15274, 16'd10993, 16'd29147, 16'd26631, 16'd42920, 16'd25260, 16'd50728, 16'd57943, 16'd61597, 16'd42406}; // indx = 2055
    #10;
    addra = 32'd65792;
    dina = {96'd0, 16'd9262, 16'd871, 16'd47417, 16'd54888, 16'd50447, 16'd43063, 16'd46443, 16'd23263, 16'd33317, 16'd23649}; // indx = 2056
    #10;
    addra = 32'd65824;
    dina = {96'd0, 16'd3035, 16'd8528, 16'd14499, 16'd200, 16'd22648, 16'd3539, 16'd60689, 16'd62175, 16'd225, 16'd17961}; // indx = 2057
    #10;
    addra = 32'd65856;
    dina = {96'd0, 16'd56762, 16'd36465, 16'd34379, 16'd53383, 16'd49847, 16'd56400, 16'd53360, 16'd58534, 16'd37379, 16'd52888}; // indx = 2058
    #10;
    addra = 32'd65888;
    dina = {96'd0, 16'd53473, 16'd52446, 16'd24126, 16'd2529, 16'd63945, 16'd64584, 16'd60237, 16'd15714, 16'd6047, 16'd23535}; // indx = 2059
    #10;
    addra = 32'd65920;
    dina = {96'd0, 16'd17409, 16'd27681, 16'd64543, 16'd10272, 16'd26010, 16'd44950, 16'd45866, 16'd39754, 16'd18345, 16'd9875}; // indx = 2060
    #10;
    addra = 32'd65952;
    dina = {96'd0, 16'd8772, 16'd9470, 16'd17505, 16'd37354, 16'd58523, 16'd54832, 16'd12756, 16'd41875, 16'd12020, 16'd8783}; // indx = 2061
    #10;
    addra = 32'd65984;
    dina = {96'd0, 16'd43557, 16'd64692, 16'd2195, 16'd39347, 16'd29214, 16'd14432, 16'd32987, 16'd5897, 16'd59141, 16'd24343}; // indx = 2062
    #10;
    addra = 32'd66016;
    dina = {96'd0, 16'd384, 16'd12969, 16'd22439, 16'd11286, 16'd24854, 16'd8880, 16'd17212, 16'd36278, 16'd58862, 16'd32366}; // indx = 2063
    #10;
    addra = 32'd66048;
    dina = {96'd0, 16'd16114, 16'd10490, 16'd20115, 16'd52191, 16'd38081, 16'd43644, 16'd19482, 16'd15879, 16'd38612, 16'd30055}; // indx = 2064
    #10;
    addra = 32'd66080;
    dina = {96'd0, 16'd25513, 16'd16957, 16'd36192, 16'd4794, 16'd46841, 16'd28911, 16'd39757, 16'd32833, 16'd50170, 16'd51678}; // indx = 2065
    #10;
    addra = 32'd66112;
    dina = {96'd0, 16'd49126, 16'd42319, 16'd10388, 16'd36292, 16'd57398, 16'd56330, 16'd13127, 16'd25424, 16'd18595, 16'd5577}; // indx = 2066
    #10;
    addra = 32'd66144;
    dina = {96'd0, 16'd11075, 16'd63026, 16'd64008, 16'd12763, 16'd3760, 16'd48249, 16'd14522, 16'd15939, 16'd20023, 16'd19629}; // indx = 2067
    #10;
    addra = 32'd66176;
    dina = {96'd0, 16'd24613, 16'd48296, 16'd30933, 16'd21293, 16'd2836, 16'd56093, 16'd18734, 16'd61451, 16'd27607, 16'd28698}; // indx = 2068
    #10;
    addra = 32'd66208;
    dina = {96'd0, 16'd16448, 16'd1059, 16'd8245, 16'd53885, 16'd63045, 16'd5043, 16'd37874, 16'd48361, 16'd48260, 16'd40374}; // indx = 2069
    #10;
    addra = 32'd66240;
    dina = {96'd0, 16'd4279, 16'd2752, 16'd61721, 16'd57603, 16'd12885, 16'd54535, 16'd27226, 16'd45131, 16'd16427, 16'd9028}; // indx = 2070
    #10;
    addra = 32'd66272;
    dina = {96'd0, 16'd44337, 16'd50176, 16'd22973, 16'd21883, 16'd61811, 16'd36736, 16'd37507, 16'd42916, 16'd64416, 16'd17510}; // indx = 2071
    #10;
    addra = 32'd66304;
    dina = {96'd0, 16'd31794, 16'd43613, 16'd6491, 16'd7824, 16'd38542, 16'd39786, 16'd56310, 16'd40781, 16'd28704, 16'd60246}; // indx = 2072
    #10;
    addra = 32'd66336;
    dina = {96'd0, 16'd35830, 16'd43189, 16'd64715, 16'd21630, 16'd26231, 16'd36840, 16'd65487, 16'd63013, 16'd15620, 16'd17466}; // indx = 2073
    #10;
    addra = 32'd66368;
    dina = {96'd0, 16'd47091, 16'd26463, 16'd4842, 16'd16430, 16'd29346, 16'd52970, 16'd11588, 16'd14841, 16'd25719, 16'd16208}; // indx = 2074
    #10;
    addra = 32'd66400;
    dina = {96'd0, 16'd33593, 16'd15055, 16'd59710, 16'd11457, 16'd10978, 16'd26674, 16'd57420, 16'd37628, 16'd1624, 16'd11997}; // indx = 2075
    #10;
    addra = 32'd66432;
    dina = {96'd0, 16'd16436, 16'd11750, 16'd14945, 16'd44465, 16'd14197, 16'd48668, 16'd25380, 16'd28301, 16'd20039, 16'd46128}; // indx = 2076
    #10;
    addra = 32'd66464;
    dina = {96'd0, 16'd7305, 16'd3432, 16'd63253, 16'd57291, 16'd63012, 16'd41079, 16'd35639, 16'd59625, 16'd42327, 16'd44358}; // indx = 2077
    #10;
    addra = 32'd66496;
    dina = {96'd0, 16'd14101, 16'd59694, 16'd34927, 16'd45322, 16'd33724, 16'd65319, 16'd23439, 16'd35937, 16'd54696, 16'd2756}; // indx = 2078
    #10;
    addra = 32'd66528;
    dina = {96'd0, 16'd10755, 16'd1844, 16'd13163, 16'd18122, 16'd17093, 16'd18596, 16'd27057, 16'd54382, 16'd47750, 16'd14922}; // indx = 2079
    #10;
    addra = 32'd66560;
    dina = {96'd0, 16'd49062, 16'd48454, 16'd52760, 16'd54069, 16'd64413, 16'd25524, 16'd50846, 16'd49279, 16'd43791, 16'd60284}; // indx = 2080
    #10;
    addra = 32'd66592;
    dina = {96'd0, 16'd56027, 16'd51161, 16'd10249, 16'd14145, 16'd57193, 16'd31968, 16'd32739, 16'd54574, 16'd7098, 16'd34058}; // indx = 2081
    #10;
    addra = 32'd66624;
    dina = {96'd0, 16'd63870, 16'd45614, 16'd37225, 16'd54375, 16'd6201, 16'd36743, 16'd41175, 16'd63533, 16'd65325, 16'd28305}; // indx = 2082
    #10;
    addra = 32'd66656;
    dina = {96'd0, 16'd39197, 16'd5877, 16'd57094, 16'd26827, 16'd19780, 16'd42391, 16'd3199, 16'd65128, 16'd17514, 16'd20536}; // indx = 2083
    #10;
    addra = 32'd66688;
    dina = {96'd0, 16'd13178, 16'd6002, 16'd37062, 16'd37409, 16'd2089, 16'd19384, 16'd36612, 16'd27269, 16'd49857, 16'd23859}; // indx = 2084
    #10;
    addra = 32'd66720;
    dina = {96'd0, 16'd40793, 16'd13070, 16'd58254, 16'd4588, 16'd9916, 16'd55118, 16'd29940, 16'd24849, 16'd7318, 16'd30078}; // indx = 2085
    #10;
    addra = 32'd66752;
    dina = {96'd0, 16'd36117, 16'd13025, 16'd17565, 16'd25253, 16'd8752, 16'd50683, 16'd29456, 16'd5625, 16'd24722, 16'd13978}; // indx = 2086
    #10;
    addra = 32'd66784;
    dina = {96'd0, 16'd47515, 16'd3032, 16'd5416, 16'd49643, 16'd3860, 16'd24817, 16'd34966, 16'd46555, 16'd34594, 16'd55878}; // indx = 2087
    #10;
    addra = 32'd66816;
    dina = {96'd0, 16'd19035, 16'd31442, 16'd50227, 16'd36511, 16'd13165, 16'd29026, 16'd26317, 16'd18644, 16'd39962, 16'd35768}; // indx = 2088
    #10;
    addra = 32'd66848;
    dina = {96'd0, 16'd15435, 16'd30653, 16'd11803, 16'd36448, 16'd36782, 16'd46791, 16'd22306, 16'd52382, 16'd54720, 16'd42942}; // indx = 2089
    #10;
    addra = 32'd66880;
    dina = {96'd0, 16'd23456, 16'd25530, 16'd5954, 16'd36771, 16'd62890, 16'd27835, 16'd32242, 16'd19416, 16'd25273, 16'd24785}; // indx = 2090
    #10;
    addra = 32'd66912;
    dina = {96'd0, 16'd53916, 16'd17937, 16'd32828, 16'd5275, 16'd29875, 16'd39023, 16'd17347, 16'd21858, 16'd33331, 16'd18109}; // indx = 2091
    #10;
    addra = 32'd66944;
    dina = {96'd0, 16'd19025, 16'd16786, 16'd26421, 16'd34047, 16'd23428, 16'd54547, 16'd48770, 16'd28168, 16'd12612, 16'd2350}; // indx = 2092
    #10;
    addra = 32'd66976;
    dina = {96'd0, 16'd35896, 16'd21878, 16'd49400, 16'd17268, 16'd25094, 16'd64087, 16'd30975, 16'd24305, 16'd53228, 16'd24439}; // indx = 2093
    #10;
    addra = 32'd67008;
    dina = {96'd0, 16'd45768, 16'd36925, 16'd32005, 16'd15937, 16'd37919, 16'd34184, 16'd53252, 16'd4952, 16'd36887, 16'd13406}; // indx = 2094
    #10;
    addra = 32'd67040;
    dina = {96'd0, 16'd64158, 16'd49156, 16'd9183, 16'd23146, 16'd35549, 16'd42226, 16'd2973, 16'd5378, 16'd61745, 16'd62065}; // indx = 2095
    #10;
    addra = 32'd67072;
    dina = {96'd0, 16'd8657, 16'd27775, 16'd58174, 16'd2493, 16'd5880, 16'd31270, 16'd59904, 16'd713, 16'd49119, 16'd25167}; // indx = 2096
    #10;
    addra = 32'd67104;
    dina = {96'd0, 16'd65371, 16'd62812, 16'd46192, 16'd61611, 16'd36722, 16'd10591, 16'd63466, 16'd48375, 16'd32378, 16'd17524}; // indx = 2097
    #10;
    addra = 32'd67136;
    dina = {96'd0, 16'd35610, 16'd23641, 16'd25022, 16'd21248, 16'd29238, 16'd59242, 16'd14680, 16'd30511, 16'd58784, 16'd63469}; // indx = 2098
    #10;
    addra = 32'd67168;
    dina = {96'd0, 16'd1368, 16'd1226, 16'd36390, 16'd2882, 16'd30030, 16'd42440, 16'd49097, 16'd40371, 16'd21603, 16'd57098}; // indx = 2099
    #10;
    addra = 32'd67200;
    dina = {96'd0, 16'd62089, 16'd63279, 16'd58789, 16'd8325, 16'd42718, 16'd21432, 16'd35799, 16'd15502, 16'd45376, 16'd3652}; // indx = 2100
    #10;
    addra = 32'd67232;
    dina = {96'd0, 16'd59448, 16'd37236, 16'd13627, 16'd16492, 16'd57937, 16'd33986, 16'd41120, 16'd2823, 16'd9444, 16'd13062}; // indx = 2101
    #10;
    addra = 32'd67264;
    dina = {96'd0, 16'd55110, 16'd16605, 16'd48464, 16'd801, 16'd45800, 16'd39174, 16'd42119, 16'd10461, 16'd16043, 16'd8653}; // indx = 2102
    #10;
    addra = 32'd67296;
    dina = {96'd0, 16'd36556, 16'd48591, 16'd34685, 16'd65085, 16'd42751, 16'd38194, 16'd3363, 16'd61130, 16'd32358, 16'd48540}; // indx = 2103
    #10;
    addra = 32'd67328;
    dina = {96'd0, 16'd8243, 16'd5981, 16'd28728, 16'd57192, 16'd40647, 16'd5116, 16'd64016, 16'd37673, 16'd18475, 16'd38929}; // indx = 2104
    #10;
    addra = 32'd67360;
    dina = {96'd0, 16'd258, 16'd27933, 16'd13487, 16'd14236, 16'd21290, 16'd48450, 16'd16595, 16'd38929, 16'd39700, 16'd65514}; // indx = 2105
    #10;
    addra = 32'd67392;
    dina = {96'd0, 16'd21469, 16'd28551, 16'd58676, 16'd56321, 16'd20105, 16'd1944, 16'd8766, 16'd12530, 16'd59500, 16'd64902}; // indx = 2106
    #10;
    addra = 32'd67424;
    dina = {96'd0, 16'd24776, 16'd31611, 16'd57339, 16'd40902, 16'd22356, 16'd15213, 16'd36575, 16'd31449, 16'd57772, 16'd36178}; // indx = 2107
    #10;
    addra = 32'd67456;
    dina = {96'd0, 16'd57028, 16'd27948, 16'd37938, 16'd16827, 16'd41142, 16'd36329, 16'd62161, 16'd8668, 16'd45112, 16'd4247}; // indx = 2108
    #10;
    addra = 32'd67488;
    dina = {96'd0, 16'd7228, 16'd45902, 16'd53273, 16'd15307, 16'd65371, 16'd43115, 16'd33931, 16'd23743, 16'd7240, 16'd54942}; // indx = 2109
    #10;
    addra = 32'd67520;
    dina = {96'd0, 16'd53785, 16'd25670, 16'd27343, 16'd31312, 16'd1341, 16'd63895, 16'd23200, 16'd54871, 16'd21799, 16'd55483}; // indx = 2110
    #10;
    addra = 32'd67552;
    dina = {96'd0, 16'd20679, 16'd3282, 16'd62826, 16'd40215, 16'd18594, 16'd20144, 16'd6937, 16'd45121, 16'd63385, 16'd25367}; // indx = 2111
    #10;
    addra = 32'd67584;
    dina = {96'd0, 16'd11551, 16'd45584, 16'd53209, 16'd27218, 16'd19850, 16'd17994, 16'd28279, 16'd11015, 16'd3196, 16'd41147}; // indx = 2112
    #10;
    addra = 32'd67616;
    dina = {96'd0, 16'd24386, 16'd40893, 16'd27244, 16'd49393, 16'd8080, 16'd26558, 16'd41850, 16'd63640, 16'd49302, 16'd46326}; // indx = 2113
    #10;
    addra = 32'd67648;
    dina = {96'd0, 16'd33256, 16'd51415, 16'd7787, 16'd32306, 16'd57454, 16'd14610, 16'd18712, 16'd17147, 16'd49994, 16'd44588}; // indx = 2114
    #10;
    addra = 32'd67680;
    dina = {96'd0, 16'd45165, 16'd56938, 16'd925, 16'd16963, 16'd7474, 16'd27813, 16'd29926, 16'd52292, 16'd38096, 16'd156}; // indx = 2115
    #10;
    addra = 32'd67712;
    dina = {96'd0, 16'd49776, 16'd17086, 16'd25796, 16'd16690, 16'd54016, 16'd54286, 16'd10002, 16'd52089, 16'd53416, 16'd64916}; // indx = 2116
    #10;
    addra = 32'd67744;
    dina = {96'd0, 16'd62912, 16'd43344, 16'd45638, 16'd48992, 16'd42857, 16'd61291, 16'd18356, 16'd42659, 16'd63530, 16'd4758}; // indx = 2117
    #10;
    addra = 32'd67776;
    dina = {96'd0, 16'd3672, 16'd58215, 16'd49201, 16'd54992, 16'd11971, 16'd26696, 16'd39087, 16'd37473, 16'd44409, 16'd54428}; // indx = 2118
    #10;
    addra = 32'd67808;
    dina = {96'd0, 16'd54968, 16'd53040, 16'd20179, 16'd14581, 16'd14823, 16'd9179, 16'd6961, 16'd32584, 16'd29484, 16'd32588}; // indx = 2119
    #10;
    addra = 32'd67840;
    dina = {96'd0, 16'd57703, 16'd22267, 16'd2827, 16'd24499, 16'd33397, 16'd64522, 16'd32860, 16'd17078, 16'd2027, 16'd34737}; // indx = 2120
    #10;
    addra = 32'd67872;
    dina = {96'd0, 16'd59104, 16'd29333, 16'd57510, 16'd61725, 16'd37170, 16'd24123, 16'd54490, 16'd15785, 16'd21790, 16'd32510}; // indx = 2121
    #10;
    addra = 32'd67904;
    dina = {96'd0, 16'd13477, 16'd28663, 16'd7445, 16'd5326, 16'd40178, 16'd54258, 16'd33026, 16'd6501, 16'd64881, 16'd2607}; // indx = 2122
    #10;
    addra = 32'd67936;
    dina = {96'd0, 16'd2193, 16'd56146, 16'd28390, 16'd48022, 16'd37652, 16'd48331, 16'd56875, 16'd42166, 16'd60777, 16'd46618}; // indx = 2123
    #10;
    addra = 32'd67968;
    dina = {96'd0, 16'd9284, 16'd15328, 16'd8603, 16'd63234, 16'd2220, 16'd49813, 16'd25867, 16'd12476, 16'd54478, 16'd9862}; // indx = 2124
    #10;
    addra = 32'd68000;
    dina = {96'd0, 16'd5605, 16'd45117, 16'd1745, 16'd20050, 16'd34296, 16'd63958, 16'd23467, 16'd37815, 16'd64137, 16'd28113}; // indx = 2125
    #10;
    addra = 32'd68032;
    dina = {96'd0, 16'd36042, 16'd21278, 16'd16167, 16'd12177, 16'd43331, 16'd15665, 16'd31347, 16'd33409, 16'd63090, 16'd48536}; // indx = 2126
    #10;
    addra = 32'd68064;
    dina = {96'd0, 16'd39034, 16'd65426, 16'd48856, 16'd40835, 16'd34250, 16'd5481, 16'd33326, 16'd4526, 16'd12999, 16'd57118}; // indx = 2127
    #10;
    addra = 32'd68096;
    dina = {96'd0, 16'd20703, 16'd39413, 16'd47385, 16'd40498, 16'd62829, 16'd7601, 16'd13423, 16'd442, 16'd32137, 16'd29222}; // indx = 2128
    #10;
    addra = 32'd68128;
    dina = {96'd0, 16'd45275, 16'd7682, 16'd20294, 16'd12743, 16'd62711, 16'd1831, 16'd11247, 16'd63550, 16'd4406, 16'd35975}; // indx = 2129
    #10;
    addra = 32'd68160;
    dina = {96'd0, 16'd6149, 16'd19890, 16'd8960, 16'd24983, 16'd52007, 16'd19735, 16'd6012, 16'd30816, 16'd31794, 16'd57154}; // indx = 2130
    #10;
    addra = 32'd68192;
    dina = {96'd0, 16'd54653, 16'd45477, 16'd27694, 16'd47183, 16'd28216, 16'd22598, 16'd13025, 16'd19101, 16'd50784, 16'd44785}; // indx = 2131
    #10;
    addra = 32'd68224;
    dina = {96'd0, 16'd55429, 16'd50460, 16'd51936, 16'd24043, 16'd20117, 16'd36975, 16'd64162, 16'd22167, 16'd39840, 16'd51670}; // indx = 2132
    #10;
    addra = 32'd68256;
    dina = {96'd0, 16'd23015, 16'd802, 16'd17179, 16'd59443, 16'd1370, 16'd54631, 16'd37562, 16'd9415, 16'd23533, 16'd6890}; // indx = 2133
    #10;
    addra = 32'd68288;
    dina = {96'd0, 16'd1717, 16'd50898, 16'd24280, 16'd8090, 16'd57779, 16'd25136, 16'd48467, 16'd58222, 16'd33941, 16'd61347}; // indx = 2134
    #10;
    addra = 32'd68320;
    dina = {96'd0, 16'd62022, 16'd47657, 16'd48103, 16'd23072, 16'd46692, 16'd18231, 16'd51110, 16'd54762, 16'd48809, 16'd38812}; // indx = 2135
    #10;
    addra = 32'd68352;
    dina = {96'd0, 16'd8878, 16'd51741, 16'd27536, 16'd14373, 16'd5921, 16'd44159, 16'd5067, 16'd5569, 16'd44313, 16'd5587}; // indx = 2136
    #10;
    addra = 32'd68384;
    dina = {96'd0, 16'd6886, 16'd54328, 16'd61780, 16'd50466, 16'd18808, 16'd37152, 16'd6265, 16'd8232, 16'd29587, 16'd8250}; // indx = 2137
    #10;
    addra = 32'd68416;
    dina = {96'd0, 16'd8487, 16'd61968, 16'd19488, 16'd8716, 16'd46810, 16'd20742, 16'd60472, 16'd25475, 16'd52055, 16'd61761}; // indx = 2138
    #10;
    addra = 32'd68448;
    dina = {96'd0, 16'd266, 16'd42557, 16'd5570, 16'd3603, 16'd38468, 16'd44003, 16'd15711, 16'd50909, 16'd56290, 16'd32499}; // indx = 2139
    #10;
    addra = 32'd68480;
    dina = {96'd0, 16'd60317, 16'd55192, 16'd45131, 16'd48218, 16'd31193, 16'd30013, 16'd5908, 16'd23649, 16'd54143, 16'd24498}; // indx = 2140
    #10;
    addra = 32'd68512;
    dina = {96'd0, 16'd23818, 16'd18544, 16'd37314, 16'd57428, 16'd37328, 16'd58438, 16'd10897, 16'd1368, 16'd3500, 16'd51598}; // indx = 2141
    #10;
    addra = 32'd68544;
    dina = {96'd0, 16'd38448, 16'd44617, 16'd26444, 16'd59731, 16'd6461, 16'd59606, 16'd24562, 16'd13031, 16'd17066, 16'd63538}; // indx = 2142
    #10;
    addra = 32'd68576;
    dina = {96'd0, 16'd38141, 16'd48332, 16'd13876, 16'd30250, 16'd8688, 16'd53403, 16'd57764, 16'd47585, 16'd32968, 16'd5656}; // indx = 2143
    #10;
    addra = 32'd68608;
    dina = {96'd0, 16'd49028, 16'd34449, 16'd2349, 16'd12122, 16'd36326, 16'd13351, 16'd22465, 16'd43756, 16'd29948, 16'd48987}; // indx = 2144
    #10;
    addra = 32'd68640;
    dina = {96'd0, 16'd34885, 16'd32357, 16'd24358, 16'd22838, 16'd23951, 16'd54078, 16'd5334, 16'd3544, 16'd32118, 16'd36042}; // indx = 2145
    #10;
    addra = 32'd68672;
    dina = {96'd0, 16'd56096, 16'd38557, 16'd2846, 16'd26823, 16'd64253, 16'd53523, 16'd27670, 16'd15838, 16'd63534, 16'd53321}; // indx = 2146
    #10;
    addra = 32'd68704;
    dina = {96'd0, 16'd56043, 16'd42866, 16'd14029, 16'd47620, 16'd56403, 16'd15808, 16'd3021, 16'd61219, 16'd16598, 16'd11797}; // indx = 2147
    #10;
    addra = 32'd68736;
    dina = {96'd0, 16'd10320, 16'd43610, 16'd22409, 16'd23621, 16'd45497, 16'd41585, 16'd52396, 16'd25756, 16'd53221, 16'd30249}; // indx = 2148
    #10;
    addra = 32'd68768;
    dina = {96'd0, 16'd18589, 16'd30329, 16'd40302, 16'd55996, 16'd59164, 16'd15166, 16'd3302, 16'd11168, 16'd32261, 16'd16394}; // indx = 2149
    #10;
    addra = 32'd68800;
    dina = {96'd0, 16'd64633, 16'd3476, 16'd33718, 16'd9883, 16'd6409, 16'd38616, 16'd11272, 16'd10533, 16'd20610, 16'd45833}; // indx = 2150
    #10;
    addra = 32'd68832;
    dina = {96'd0, 16'd52290, 16'd46162, 16'd7292, 16'd30571, 16'd52621, 16'd47473, 16'd8593, 16'd18934, 16'd32686, 16'd44720}; // indx = 2151
    #10;
    addra = 32'd68864;
    dina = {96'd0, 16'd4834, 16'd8110, 16'd57360, 16'd18719, 16'd22773, 16'd58371, 16'd28724, 16'd36580, 16'd7882, 16'd9832}; // indx = 2152
    #10;
    addra = 32'd68896;
    dina = {96'd0, 16'd5719, 16'd62590, 16'd64413, 16'd61893, 16'd64963, 16'd64434, 16'd11614, 16'd22787, 16'd40060, 16'd52219}; // indx = 2153
    #10;
    addra = 32'd68928;
    dina = {96'd0, 16'd19310, 16'd27232, 16'd59651, 16'd15773, 16'd23114, 16'd17917, 16'd40632, 16'd30132, 16'd15784, 16'd53672}; // indx = 2154
    #10;
    addra = 32'd68960;
    dina = {96'd0, 16'd39746, 16'd37178, 16'd50000, 16'd17357, 16'd47719, 16'd61922, 16'd55184, 16'd5079, 16'd48347, 16'd17275}; // indx = 2155
    #10;
    addra = 32'd68992;
    dina = {96'd0, 16'd60925, 16'd13, 16'd45226, 16'd28191, 16'd50116, 16'd45422, 16'd55726, 16'd64083, 16'd23626, 16'd41907}; // indx = 2156
    #10;
    addra = 32'd69024;
    dina = {96'd0, 16'd11780, 16'd56664, 16'd28181, 16'd55348, 16'd53105, 16'd35875, 16'd40674, 16'd1716, 16'd23045, 16'd26002}; // indx = 2157
    #10;
    addra = 32'd69056;
    dina = {96'd0, 16'd58347, 16'd12886, 16'd36432, 16'd62862, 16'd18573, 16'd34061, 16'd6815, 16'd45643, 16'd32144, 16'd16273}; // indx = 2158
    #10;
    addra = 32'd69088;
    dina = {96'd0, 16'd53845, 16'd38741, 16'd13542, 16'd61672, 16'd3244, 16'd16075, 16'd43449, 16'd25782, 16'd52769, 16'd21540}; // indx = 2159
    #10;
    addra = 32'd69120;
    dina = {96'd0, 16'd42704, 16'd5035, 16'd23315, 16'd225, 16'd5505, 16'd58114, 16'd38823, 16'd44045, 16'd19832, 16'd28120}; // indx = 2160
    #10;
    addra = 32'd69152;
    dina = {96'd0, 16'd45407, 16'd48529, 16'd7395, 16'd1185, 16'd44708, 16'd25132, 16'd59657, 16'd15473, 16'd37629, 16'd26523}; // indx = 2161
    #10;
    addra = 32'd69184;
    dina = {96'd0, 16'd40109, 16'd21145, 16'd22902, 16'd46805, 16'd21652, 16'd44004, 16'd18030, 16'd18670, 16'd24866, 16'd5559}; // indx = 2162
    #10;
    addra = 32'd69216;
    dina = {96'd0, 16'd1990, 16'd34754, 16'd27908, 16'd6910, 16'd36074, 16'd47795, 16'd28613, 16'd54455, 16'd43864, 16'd49211}; // indx = 2163
    #10;
    addra = 32'd69248;
    dina = {96'd0, 16'd48208, 16'd38422, 16'd23723, 16'd51200, 16'd4413, 16'd34236, 16'd46606, 16'd48644, 16'd63512, 16'd1}; // indx = 2164
    #10;
    addra = 32'd69280;
    dina = {96'd0, 16'd55053, 16'd26298, 16'd54886, 16'd1938, 16'd29347, 16'd36965, 16'd2220, 16'd41404, 16'd32078, 16'd19172}; // indx = 2165
    #10;
    addra = 32'd69312;
    dina = {96'd0, 16'd37383, 16'd53316, 16'd64573, 16'd41860, 16'd61263, 16'd4902, 16'd56331, 16'd13347, 16'd38119, 16'd23460}; // indx = 2166
    #10;
    addra = 32'd69344;
    dina = {96'd0, 16'd47695, 16'd46377, 16'd33725, 16'd33563, 16'd12774, 16'd12115, 16'd21682, 16'd3736, 16'd58274, 16'd16867}; // indx = 2167
    #10;
    addra = 32'd69376;
    dina = {96'd0, 16'd36822, 16'd18145, 16'd1919, 16'd12049, 16'd50137, 16'd50632, 16'd46223, 16'd63775, 16'd54658, 16'd57545}; // indx = 2168
    #10;
    addra = 32'd69408;
    dina = {96'd0, 16'd36096, 16'd11058, 16'd23238, 16'd23883, 16'd36425, 16'd50383, 16'd49654, 16'd62399, 16'd17996, 16'd7820}; // indx = 2169
    #10;
    addra = 32'd69440;
    dina = {96'd0, 16'd7335, 16'd53022, 16'd26250, 16'd43920, 16'd29032, 16'd1456, 16'd10886, 16'd37316, 16'd45977, 16'd42867}; // indx = 2170
    #10;
    addra = 32'd69472;
    dina = {96'd0, 16'd5299, 16'd29728, 16'd56453, 16'd23949, 16'd15653, 16'd54932, 16'd11323, 16'd5628, 16'd37508, 16'd35202}; // indx = 2171
    #10;
    addra = 32'd69504;
    dina = {96'd0, 16'd39311, 16'd18915, 16'd50977, 16'd33119, 16'd53064, 16'd53180, 16'd37657, 16'd44469, 16'd25393, 16'd46734}; // indx = 2172
    #10;
    addra = 32'd69536;
    dina = {96'd0, 16'd8687, 16'd29950, 16'd26751, 16'd17275, 16'd21489, 16'd55143, 16'd29440, 16'd28819, 16'd36756, 16'd45913}; // indx = 2173
    #10;
    addra = 32'd69568;
    dina = {96'd0, 16'd49706, 16'd64504, 16'd63541, 16'd49171, 16'd6859, 16'd43484, 16'd60588, 16'd53312, 16'd56876, 16'd60861}; // indx = 2174
    #10;
    addra = 32'd69600;
    dina = {96'd0, 16'd54354, 16'd18521, 16'd14032, 16'd34780, 16'd57388, 16'd30980, 16'd32172, 16'd11699, 16'd26753, 16'd875}; // indx = 2175
    #10;
    addra = 32'd69632;
    dina = {96'd0, 16'd31415, 16'd24571, 16'd39674, 16'd27021, 16'd52904, 16'd19270, 16'd58870, 16'd44474, 16'd14998, 16'd21158}; // indx = 2176
    #10;
    addra = 32'd69664;
    dina = {96'd0, 16'd1674, 16'd24333, 16'd58785, 16'd60066, 16'd32466, 16'd22657, 16'd50077, 16'd63190, 16'd10448, 16'd13226}; // indx = 2177
    #10;
    addra = 32'd69696;
    dina = {96'd0, 16'd65450, 16'd38554, 16'd60029, 16'd45863, 16'd51079, 16'd12093, 16'd47053, 16'd31014, 16'd30433, 16'd24785}; // indx = 2178
    #10;
    addra = 32'd69728;
    dina = {96'd0, 16'd48783, 16'd43226, 16'd41531, 16'd50957, 16'd43152, 16'd21130, 16'd28327, 16'd43482, 16'd26856, 16'd42566}; // indx = 2179
    #10;
    addra = 32'd69760;
    dina = {96'd0, 16'd22334, 16'd11054, 16'd33278, 16'd54396, 16'd54451, 16'd522, 16'd45417, 16'd15353, 16'd7415, 16'd40266}; // indx = 2180
    #10;
    addra = 32'd69792;
    dina = {96'd0, 16'd2927, 16'd28063, 16'd45026, 16'd19479, 16'd44605, 16'd27168, 16'd16021, 16'd47383, 16'd40435, 16'd60596}; // indx = 2181
    #10;
    addra = 32'd69824;
    dina = {96'd0, 16'd47063, 16'd16377, 16'd33932, 16'd38509, 16'd13744, 16'd31880, 16'd5585, 16'd24179, 16'd27141, 16'd32647}; // indx = 2182
    #10;
    addra = 32'd69856;
    dina = {96'd0, 16'd64252, 16'd38747, 16'd58097, 16'd20223, 16'd27520, 16'd34833, 16'd20874, 16'd60242, 16'd31687, 16'd41509}; // indx = 2183
    #10;
    addra = 32'd69888;
    dina = {96'd0, 16'd15201, 16'd51758, 16'd46835, 16'd57668, 16'd8472, 16'd34845, 16'd45004, 16'd12805, 16'd58306, 16'd18431}; // indx = 2184
    #10;
    addra = 32'd69920;
    dina = {96'd0, 16'd24967, 16'd8684, 16'd4103, 16'd65150, 16'd36083, 16'd35166, 16'd31607, 16'd60784, 16'd5773, 16'd36513}; // indx = 2185
    #10;
    addra = 32'd69952;
    dina = {96'd0, 16'd12118, 16'd45337, 16'd22826, 16'd38794, 16'd38964, 16'd15052, 16'd21879, 16'd10459, 16'd37713, 16'd62547}; // indx = 2186
    #10;
    addra = 32'd69984;
    dina = {96'd0, 16'd56398, 16'd27094, 16'd13011, 16'd21879, 16'd53311, 16'd28484, 16'd8498, 16'd9513, 16'd30727, 16'd13221}; // indx = 2187
    #10;
    addra = 32'd70016;
    dina = {96'd0, 16'd24160, 16'd55297, 16'd29498, 16'd16879, 16'd2835, 16'd28620, 16'd62964, 16'd46299, 16'd47850, 16'd3064}; // indx = 2188
    #10;
    addra = 32'd70048;
    dina = {96'd0, 16'd60187, 16'd9896, 16'd29036, 16'd40387, 16'd21577, 16'd40319, 16'd60735, 16'd7089, 16'd45038, 16'd55630}; // indx = 2189
    #10;
    addra = 32'd70080;
    dina = {96'd0, 16'd48865, 16'd65390, 16'd48208, 16'd41714, 16'd20495, 16'd17845, 16'd7896, 16'd42431, 16'd20197, 16'd56099}; // indx = 2190
    #10;
    addra = 32'd70112;
    dina = {96'd0, 16'd58679, 16'd47455, 16'd53718, 16'd52545, 16'd53746, 16'd19545, 16'd21224, 16'd44326, 16'd15372, 16'd8587}; // indx = 2191
    #10;
    addra = 32'd70144;
    dina = {96'd0, 16'd23198, 16'd52766, 16'd29786, 16'd14525, 16'd40963, 16'd18809, 16'd25035, 16'd37893, 16'd29248, 16'd21627}; // indx = 2192
    #10;
    addra = 32'd70176;
    dina = {96'd0, 16'd61845, 16'd29348, 16'd8360, 16'd32646, 16'd23007, 16'd5953, 16'd64218, 16'd13169, 16'd42306, 16'd29140}; // indx = 2193
    #10;
    addra = 32'd70208;
    dina = {96'd0, 16'd44657, 16'd12987, 16'd23865, 16'd59777, 16'd56223, 16'd4709, 16'd23701, 16'd37641, 16'd47726, 16'd45400}; // indx = 2194
    #10;
    addra = 32'd70240;
    dina = {96'd0, 16'd18042, 16'd34537, 16'd51325, 16'd4291, 16'd11568, 16'd3779, 16'd17160, 16'd20059, 16'd14024, 16'd41471}; // indx = 2195
    #10;
    addra = 32'd70272;
    dina = {96'd0, 16'd61683, 16'd46314, 16'd61826, 16'd14556, 16'd12445, 16'd23102, 16'd53068, 16'd54222, 16'd29590, 16'd24130}; // indx = 2196
    #10;
    addra = 32'd70304;
    dina = {96'd0, 16'd54159, 16'd54980, 16'd40529, 16'd16375, 16'd7287, 16'd46003, 16'd52590, 16'd43540, 16'd53384, 16'd13837}; // indx = 2197
    #10;
    addra = 32'd70336;
    dina = {96'd0, 16'd6979, 16'd34451, 16'd58424, 16'd9120, 16'd2053, 16'd29322, 16'd38075, 16'd25515, 16'd42838, 16'd13008}; // indx = 2198
    #10;
    addra = 32'd70368;
    dina = {96'd0, 16'd48189, 16'd9970, 16'd41355, 16'd5561, 16'd1131, 16'd14776, 16'd57794, 16'd56680, 16'd19007, 16'd49045}; // indx = 2199
    #10;
    addra = 32'd70400;
    dina = {96'd0, 16'd15792, 16'd34211, 16'd9078, 16'd13967, 16'd45947, 16'd60478, 16'd10606, 16'd51786, 16'd14226, 16'd33167}; // indx = 2200
    #10;
    addra = 32'd70432;
    dina = {96'd0, 16'd61918, 16'd42576, 16'd49797, 16'd3932, 16'd21874, 16'd53692, 16'd49984, 16'd51535, 16'd60467, 16'd46646}; // indx = 2201
    #10;
    addra = 32'd70464;
    dina = {96'd0, 16'd1270, 16'd42616, 16'd58549, 16'd11763, 16'd32294, 16'd41755, 16'd24103, 16'd23052, 16'd30548, 16'd41042}; // indx = 2202
    #10;
    addra = 32'd70496;
    dina = {96'd0, 16'd32164, 16'd46680, 16'd22982, 16'd63025, 16'd48591, 16'd26593, 16'd13037, 16'd438, 16'd53091, 16'd34285}; // indx = 2203
    #10;
    addra = 32'd70528;
    dina = {96'd0, 16'd3620, 16'd36912, 16'd62074, 16'd38602, 16'd36278, 16'd62542, 16'd34002, 16'd39913, 16'd5617, 16'd24830}; // indx = 2204
    #10;
    addra = 32'd70560;
    dina = {96'd0, 16'd27084, 16'd51792, 16'd56703, 16'd46444, 16'd7892, 16'd22149, 16'd63325, 16'd46202, 16'd38382, 16'd36302}; // indx = 2205
    #10;
    addra = 32'd70592;
    dina = {96'd0, 16'd45723, 16'd32201, 16'd53591, 16'd28946, 16'd20101, 16'd16902, 16'd26401, 16'd52248, 16'd5679, 16'd49624}; // indx = 2206
    #10;
    addra = 32'd70624;
    dina = {96'd0, 16'd52453, 16'd33314, 16'd34703, 16'd36629, 16'd31153, 16'd18874, 16'd26682, 16'd45280, 16'd37304, 16'd34513}; // indx = 2207
    #10;
    addra = 32'd70656;
    dina = {96'd0, 16'd22362, 16'd60711, 16'd54349, 16'd14753, 16'd56894, 16'd35459, 16'd34911, 16'd49210, 16'd10250, 16'd14209}; // indx = 2208
    #10;
    addra = 32'd70688;
    dina = {96'd0, 16'd7607, 16'd14141, 16'd44395, 16'd13842, 16'd18349, 16'd37222, 16'd14000, 16'd62906, 16'd48723, 16'd38529}; // indx = 2209
    #10;
    addra = 32'd70720;
    dina = {96'd0, 16'd40741, 16'd15674, 16'd15642, 16'd49799, 16'd41488, 16'd8261, 16'd51500, 16'd13606, 16'd54883, 16'd32561}; // indx = 2210
    #10;
    addra = 32'd70752;
    dina = {96'd0, 16'd39061, 16'd59035, 16'd20958, 16'd40354, 16'd41750, 16'd1776, 16'd60584, 16'd25821, 16'd24302, 16'd46168}; // indx = 2211
    #10;
    addra = 32'd70784;
    dina = {96'd0, 16'd63288, 16'd15450, 16'd53665, 16'd26260, 16'd29738, 16'd32220, 16'd54701, 16'd7448, 16'd61790, 16'd4416}; // indx = 2212
    #10;
    addra = 32'd70816;
    dina = {96'd0, 16'd39676, 16'd35802, 16'd49607, 16'd57524, 16'd40188, 16'd55384, 16'd24591, 16'd7397, 16'd7642, 16'd7931}; // indx = 2213
    #10;
    addra = 32'd70848;
    dina = {96'd0, 16'd50916, 16'd36172, 16'd36447, 16'd63564, 16'd53298, 16'd9131, 16'd3494, 16'd4592, 16'd14813, 16'd50465}; // indx = 2214
    #10;
    addra = 32'd70880;
    dina = {96'd0, 16'd21886, 16'd15170, 16'd39651, 16'd45747, 16'd25282, 16'd63785, 16'd64499, 16'd841, 16'd63531, 16'd61842}; // indx = 2215
    #10;
    addra = 32'd70912;
    dina = {96'd0, 16'd50553, 16'd62633, 16'd31313, 16'd30227, 16'd59752, 16'd19688, 16'd10402, 16'd62120, 16'd60051, 16'd36091}; // indx = 2216
    #10;
    addra = 32'd70944;
    dina = {96'd0, 16'd47019, 16'd11310, 16'd65433, 16'd30807, 16'd35943, 16'd58985, 16'd44606, 16'd808, 16'd49834, 16'd54852}; // indx = 2217
    #10;
    addra = 32'd70976;
    dina = {96'd0, 16'd29109, 16'd54030, 16'd59172, 16'd33458, 16'd62133, 16'd10, 16'd64049, 16'd63501, 16'd14093, 16'd20559}; // indx = 2218
    #10;
    addra = 32'd71008;
    dina = {96'd0, 16'd35489, 16'd20945, 16'd60833, 16'd11883, 16'd11620, 16'd9040, 16'd64945, 16'd6934, 16'd61257, 16'd40942}; // indx = 2219
    #10;
    addra = 32'd71040;
    dina = {96'd0, 16'd50759, 16'd31138, 16'd37006, 16'd18376, 16'd12965, 16'd15858, 16'd45500, 16'd43928, 16'd11332, 16'd53354}; // indx = 2220
    #10;
    addra = 32'd71072;
    dina = {96'd0, 16'd53907, 16'd10986, 16'd57257, 16'd38761, 16'd17885, 16'd26724, 16'd39564, 16'd65360, 16'd41119, 16'd46654}; // indx = 2221
    #10;
    addra = 32'd71104;
    dina = {96'd0, 16'd56675, 16'd45295, 16'd23936, 16'd22532, 16'd20164, 16'd31324, 16'd333, 16'd315, 16'd3524, 16'd65334}; // indx = 2222
    #10;
    addra = 32'd71136;
    dina = {96'd0, 16'd14110, 16'd62030, 16'd10631, 16'd10556, 16'd50689, 16'd23742, 16'd14545, 16'd51426, 16'd44164, 16'd15114}; // indx = 2223
    #10;
    addra = 32'd71168;
    dina = {96'd0, 16'd17442, 16'd49003, 16'd52886, 16'd21902, 16'd38885, 16'd45215, 16'd10147, 16'd2941, 16'd37155, 16'd12987}; // indx = 2224
    #10;
    addra = 32'd71200;
    dina = {96'd0, 16'd24423, 16'd41066, 16'd54583, 16'd41864, 16'd17199, 16'd56725, 16'd18713, 16'd13534, 16'd16624, 16'd55703}; // indx = 2225
    #10;
    addra = 32'd71232;
    dina = {96'd0, 16'd1791, 16'd46867, 16'd47059, 16'd45634, 16'd23294, 16'd40809, 16'd39777, 16'd26265, 16'd44744, 16'd7784}; // indx = 2226
    #10;
    addra = 32'd71264;
    dina = {96'd0, 16'd13704, 16'd35588, 16'd25929, 16'd57172, 16'd58743, 16'd15582, 16'd42981, 16'd3050, 16'd3967, 16'd5590}; // indx = 2227
    #10;
    addra = 32'd71296;
    dina = {96'd0, 16'd62602, 16'd479, 16'd4391, 16'd31925, 16'd5738, 16'd18801, 16'd65074, 16'd8156, 16'd60822, 16'd51374}; // indx = 2228
    #10;
    addra = 32'd71328;
    dina = {96'd0, 16'd10652, 16'd1220, 16'd34506, 16'd20763, 16'd61047, 16'd30689, 16'd59307, 16'd47710, 16'd13512, 16'd14976}; // indx = 2229
    #10;
    addra = 32'd71360;
    dina = {96'd0, 16'd3121, 16'd6011, 16'd46381, 16'd9350, 16'd40789, 16'd59989, 16'd12316, 16'd29988, 16'd6140, 16'd19753}; // indx = 2230
    #10;
    addra = 32'd71392;
    dina = {96'd0, 16'd60758, 16'd31428, 16'd63028, 16'd26400, 16'd46231, 16'd30360, 16'd21214, 16'd53892, 16'd18223, 16'd53677}; // indx = 2231
    #10;
    addra = 32'd71424;
    dina = {96'd0, 16'd14161, 16'd38506, 16'd25471, 16'd47649, 16'd53787, 16'd34048, 16'd48877, 16'd34621, 16'd12607, 16'd29487}; // indx = 2232
    #10;
    addra = 32'd71456;
    dina = {96'd0, 16'd52166, 16'd20924, 16'd22839, 16'd54988, 16'd29143, 16'd49854, 16'd27279, 16'd14527, 16'd28892, 16'd9986}; // indx = 2233
    #10;
    addra = 32'd71488;
    dina = {96'd0, 16'd19856, 16'd60853, 16'd33449, 16'd32677, 16'd62156, 16'd40753, 16'd21331, 16'd17166, 16'd36973, 16'd32224}; // indx = 2234
    #10;
    addra = 32'd71520;
    dina = {96'd0, 16'd44044, 16'd24715, 16'd25171, 16'd35270, 16'd20019, 16'd4729, 16'd59592, 16'd18706, 16'd42007, 16'd48998}; // indx = 2235
    #10;
    addra = 32'd71552;
    dina = {96'd0, 16'd35519, 16'd44565, 16'd55679, 16'd17767, 16'd38125, 16'd29772, 16'd13330, 16'd31694, 16'd58381, 16'd45372}; // indx = 2236
    #10;
    addra = 32'd71584;
    dina = {96'd0, 16'd41176, 16'd12396, 16'd46847, 16'd59614, 16'd23902, 16'd26625, 16'd55040, 16'd22263, 16'd61417, 16'd22212}; // indx = 2237
    #10;
    addra = 32'd71616;
    dina = {96'd0, 16'd10623, 16'd49769, 16'd39600, 16'd39111, 16'd12750, 16'd32787, 16'd18967, 16'd4066, 16'd64102, 16'd9363}; // indx = 2238
    #10;
    addra = 32'd71648;
    dina = {96'd0, 16'd22248, 16'd3630, 16'd33515, 16'd7494, 16'd22377, 16'd50346, 16'd17109, 16'd60065, 16'd43058, 16'd38289}; // indx = 2239
    #10;
    addra = 32'd71680;
    dina = {96'd0, 16'd44378, 16'd52729, 16'd32381, 16'd57517, 16'd23179, 16'd12137, 16'd10138, 16'd54886, 16'd37297, 16'd41093}; // indx = 2240
    #10;
    addra = 32'd71712;
    dina = {96'd0, 16'd54373, 16'd31512, 16'd26660, 16'd19603, 16'd31170, 16'd54928, 16'd50996, 16'd36487, 16'd61580, 16'd59406}; // indx = 2241
    #10;
    addra = 32'd71744;
    dina = {96'd0, 16'd50108, 16'd28831, 16'd48603, 16'd22305, 16'd36103, 16'd558, 16'd43026, 16'd19490, 16'd10219, 16'd57193}; // indx = 2242
    #10;
    addra = 32'd71776;
    dina = {96'd0, 16'd21883, 16'd55501, 16'd7437, 16'd53323, 16'd50385, 16'd51471, 16'd29985, 16'd1177, 16'd5121, 16'd30745}; // indx = 2243
    #10;
    addra = 32'd71808;
    dina = {96'd0, 16'd19121, 16'd19527, 16'd23258, 16'd6989, 16'd59362, 16'd18795, 16'd26843, 16'd11584, 16'd49099, 16'd50452}; // indx = 2244
    #10;
    addra = 32'd71840;
    dina = {96'd0, 16'd45854, 16'd29797, 16'd46480, 16'd63173, 16'd28431, 16'd10465, 16'd24721, 16'd61649, 16'd4277, 16'd24980}; // indx = 2245
    #10;
    addra = 32'd71872;
    dina = {96'd0, 16'd42420, 16'd9189, 16'd61790, 16'd2903, 16'd55289, 16'd49869, 16'd17777, 16'd58575, 16'd58486, 16'd23580}; // indx = 2246
    #10;
    addra = 32'd71904;
    dina = {96'd0, 16'd18133, 16'd47074, 16'd45997, 16'd37393, 16'd37783, 16'd6336, 16'd17626, 16'd56812, 16'd34844, 16'd28025}; // indx = 2247
    #10;
    addra = 32'd71936;
    dina = {96'd0, 16'd33264, 16'd62425, 16'd45929, 16'd23817, 16'd45661, 16'd2883, 16'd35319, 16'd56959, 16'd32297, 16'd50161}; // indx = 2248
    #10;
    addra = 32'd71968;
    dina = {96'd0, 16'd49262, 16'd43712, 16'd20862, 16'd8591, 16'd59603, 16'd2131, 16'd37682, 16'd7623, 16'd13668, 16'd24399}; // indx = 2249
    #10;
    addra = 32'd72000;
    dina = {96'd0, 16'd53772, 16'd20342, 16'd36220, 16'd729, 16'd21856, 16'd26622, 16'd36075, 16'd39167, 16'd56804, 16'd41602}; // indx = 2250
    #10;
    addra = 32'd72032;
    dina = {96'd0, 16'd43672, 16'd27694, 16'd40542, 16'd38156, 16'd50190, 16'd31871, 16'd29898, 16'd51072, 16'd2634, 16'd1945}; // indx = 2251
    #10;
    addra = 32'd72064;
    dina = {96'd0, 16'd20815, 16'd3663, 16'd42725, 16'd57737, 16'd47212, 16'd31357, 16'd3347, 16'd42492, 16'd16960, 16'd16049}; // indx = 2252
    #10;
    addra = 32'd72096;
    dina = {96'd0, 16'd50125, 16'd46882, 16'd53401, 16'd61306, 16'd61600, 16'd9519, 16'd12112, 16'd23717, 16'd56906, 16'd49156}; // indx = 2253
    #10;
    addra = 32'd72128;
    dina = {96'd0, 16'd22854, 16'd44951, 16'd43792, 16'd3591, 16'd51654, 16'd39252, 16'd46035, 16'd42927, 16'd23642, 16'd8001}; // indx = 2254
    #10;
    addra = 32'd72160;
    dina = {96'd0, 16'd5813, 16'd13272, 16'd33076, 16'd28572, 16'd58780, 16'd20392, 16'd59395, 16'd58744, 16'd20326, 16'd10999}; // indx = 2255
    #10;
    addra = 32'd72192;
    dina = {96'd0, 16'd41519, 16'd54297, 16'd47559, 16'd4160, 16'd7786, 16'd40427, 16'd53964, 16'd43814, 16'd32173, 16'd9949}; // indx = 2256
    #10;
    addra = 32'd72224;
    dina = {96'd0, 16'd14874, 16'd61186, 16'd31087, 16'd62970, 16'd12504, 16'd33515, 16'd15089, 16'd39354, 16'd45457, 16'd22469}; // indx = 2257
    #10;
    addra = 32'd72256;
    dina = {96'd0, 16'd57155, 16'd64586, 16'd23456, 16'd32406, 16'd46913, 16'd63005, 16'd9947, 16'd4995, 16'd1241, 16'd36079}; // indx = 2258
    #10;
    addra = 32'd72288;
    dina = {96'd0, 16'd33562, 16'd7581, 16'd22395, 16'd11234, 16'd10602, 16'd10903, 16'd63053, 16'd33533, 16'd15961, 16'd60659}; // indx = 2259
    #10;
    addra = 32'd72320;
    dina = {96'd0, 16'd571, 16'd7193, 16'd61434, 16'd4457, 16'd16180, 16'd21845, 16'd64219, 16'd53053, 16'd45950, 16'd40150}; // indx = 2260
    #10;
    addra = 32'd72352;
    dina = {96'd0, 16'd46827, 16'd47552, 16'd25518, 16'd6052, 16'd41625, 16'd20326, 16'd20174, 16'd13056, 16'd17141, 16'd36267}; // indx = 2261
    #10;
    addra = 32'd72384;
    dina = {96'd0, 16'd2469, 16'd59953, 16'd37896, 16'd60507, 16'd30672, 16'd23695, 16'd25685, 16'd38872, 16'd23303, 16'd59978}; // indx = 2262
    #10;
    addra = 32'd72416;
    dina = {96'd0, 16'd12624, 16'd43317, 16'd33420, 16'd39979, 16'd61956, 16'd6552, 16'd18819, 16'd23812, 16'd8440, 16'd24074}; // indx = 2263
    #10;
    addra = 32'd72448;
    dina = {96'd0, 16'd30006, 16'd41385, 16'd54114, 16'd24734, 16'd60390, 16'd26171, 16'd46867, 16'd16898, 16'd5107, 16'd8496}; // indx = 2264
    #10;
    addra = 32'd72480;
    dina = {96'd0, 16'd33814, 16'd22182, 16'd30870, 16'd53388, 16'd29019, 16'd36673, 16'd60126, 16'd17521, 16'd38518, 16'd10893}; // indx = 2265
    #10;
    addra = 32'd72512;
    dina = {96'd0, 16'd43047, 16'd45213, 16'd41010, 16'd15036, 16'd59060, 16'd57991, 16'd47969, 16'd64834, 16'd31165, 16'd13988}; // indx = 2266
    #10;
    addra = 32'd72544;
    dina = {96'd0, 16'd21893, 16'd16070, 16'd50094, 16'd49617, 16'd11707, 16'd61366, 16'd38344, 16'd65086, 16'd51956, 16'd4281}; // indx = 2267
    #10;
    addra = 32'd72576;
    dina = {96'd0, 16'd50340, 16'd54823, 16'd20716, 16'd50922, 16'd30575, 16'd59110, 16'd61579, 16'd62742, 16'd35710, 16'd33891}; // indx = 2268
    #10;
    addra = 32'd72608;
    dina = {96'd0, 16'd61901, 16'd3187, 16'd17155, 16'd60006, 16'd54022, 16'd49917, 16'd60485, 16'd7869, 16'd28933, 16'd8013}; // indx = 2269
    #10;
    addra = 32'd72640;
    dina = {96'd0, 16'd32414, 16'd27183, 16'd36051, 16'd8758, 16'd57573, 16'd48244, 16'd9149, 16'd52477, 16'd16885, 16'd9682}; // indx = 2270
    #10;
    addra = 32'd72672;
    dina = {96'd0, 16'd59471, 16'd54644, 16'd56881, 16'd36373, 16'd62796, 16'd30046, 16'd24618, 16'd63360, 16'd45120, 16'd30825}; // indx = 2271
    #10;
    addra = 32'd72704;
    dina = {96'd0, 16'd60648, 16'd52411, 16'd52243, 16'd14148, 16'd31130, 16'd47444, 16'd5008, 16'd12373, 16'd36117, 16'd13949}; // indx = 2272
    #10;
    addra = 32'd72736;
    dina = {96'd0, 16'd21680, 16'd17953, 16'd59352, 16'd60227, 16'd28483, 16'd43674, 16'd55100, 16'd32578, 16'd55746, 16'd22646}; // indx = 2273
    #10;
    addra = 32'd72768;
    dina = {96'd0, 16'd55773, 16'd59876, 16'd51217, 16'd615, 16'd44612, 16'd63123, 16'd6402, 16'd10558, 16'd27572, 16'd8009}; // indx = 2274
    #10;
    addra = 32'd72800;
    dina = {96'd0, 16'd35930, 16'd14861, 16'd50003, 16'd41692, 16'd11704, 16'd21346, 16'd25420, 16'd45600, 16'd44372, 16'd53917}; // indx = 2275
    #10;
    addra = 32'd72832;
    dina = {96'd0, 16'd57270, 16'd64222, 16'd21030, 16'd59232, 16'd7740, 16'd14945, 16'd44472, 16'd46483, 16'd64242, 16'd10401}; // indx = 2276
    #10;
    addra = 32'd72864;
    dina = {96'd0, 16'd1214, 16'd62335, 16'd60325, 16'd4457, 16'd44369, 16'd5906, 16'd51053, 16'd52381, 16'd37306, 16'd3553}; // indx = 2277
    #10;
    addra = 32'd72896;
    dina = {96'd0, 16'd49492, 16'd33673, 16'd6569, 16'd39046, 16'd49906, 16'd20477, 16'd37232, 16'd39736, 16'd37297, 16'd15280}; // indx = 2278
    #10;
    addra = 32'd72928;
    dina = {96'd0, 16'd29934, 16'd25441, 16'd57546, 16'd47454, 16'd16708, 16'd52011, 16'd45628, 16'd16013, 16'd58482, 16'd2801}; // indx = 2279
    #10;
    addra = 32'd72960;
    dina = {96'd0, 16'd52683, 16'd60648, 16'd13226, 16'd57141, 16'd48427, 16'd22404, 16'd29662, 16'd59368, 16'd46276, 16'd10466}; // indx = 2280
    #10;
    addra = 32'd72992;
    dina = {96'd0, 16'd50791, 16'd42379, 16'd32623, 16'd55946, 16'd45033, 16'd16571, 16'd48693, 16'd61562, 16'd23819, 16'd45925}; // indx = 2281
    #10;
    addra = 32'd73024;
    dina = {96'd0, 16'd125, 16'd26694, 16'd18650, 16'd25434, 16'd19956, 16'd63590, 16'd39740, 16'd40634, 16'd14054, 16'd64351}; // indx = 2282
    #10;
    addra = 32'd73056;
    dina = {96'd0, 16'd15093, 16'd6362, 16'd19737, 16'd62562, 16'd55197, 16'd62562, 16'd12257, 16'd23638, 16'd28062, 16'd16530}; // indx = 2283
    #10;
    addra = 32'd73088;
    dina = {96'd0, 16'd38302, 16'd18825, 16'd58391, 16'd15360, 16'd33929, 16'd14046, 16'd48680, 16'd22219, 16'd3927, 16'd62563}; // indx = 2284
    #10;
    addra = 32'd73120;
    dina = {96'd0, 16'd7820, 16'd23048, 16'd62538, 16'd4754, 16'd57365, 16'd46574, 16'd19914, 16'd64391, 16'd49774, 16'd11161}; // indx = 2285
    #10;
    addra = 32'd73152;
    dina = {96'd0, 16'd58972, 16'd21111, 16'd53945, 16'd25181, 16'd16679, 16'd1002, 16'd31661, 16'd3637, 16'd59845, 16'd12064}; // indx = 2286
    #10;
    addra = 32'd73184;
    dina = {96'd0, 16'd34343, 16'd30457, 16'd41094, 16'd24303, 16'd26324, 16'd63017, 16'd11070, 16'd37092, 16'd6940, 16'd34908}; // indx = 2287
    #10;
    addra = 32'd73216;
    dina = {96'd0, 16'd12556, 16'd5729, 16'd10031, 16'd32861, 16'd215, 16'd57684, 16'd46660, 16'd22937, 16'd35870, 16'd21825}; // indx = 2288
    #10;
    addra = 32'd73248;
    dina = {96'd0, 16'd8400, 16'd34749, 16'd36256, 16'd40688, 16'd54770, 16'd61410, 16'd10653, 16'd33970, 16'd3784, 16'd26865}; // indx = 2289
    #10;
    addra = 32'd73280;
    dina = {96'd0, 16'd16690, 16'd49878, 16'd9579, 16'd57487, 16'd40811, 16'd32477, 16'd18079, 16'd57841, 16'd62708, 16'd10111}; // indx = 2290
    #10;
    addra = 32'd73312;
    dina = {96'd0, 16'd2586, 16'd465, 16'd18496, 16'd59336, 16'd50978, 16'd50247, 16'd3733, 16'd30856, 16'd9762, 16'd1615}; // indx = 2291
    #10;
    addra = 32'd73344;
    dina = {96'd0, 16'd57448, 16'd31254, 16'd19049, 16'd448, 16'd4387, 16'd9719, 16'd10252, 16'd35784, 16'd38453, 16'd15846}; // indx = 2292
    #10;
    addra = 32'd73376;
    dina = {96'd0, 16'd4054, 16'd14668, 16'd3357, 16'd41721, 16'd56433, 16'd61307, 16'd4467, 16'd17860, 16'd19171, 16'd3006}; // indx = 2293
    #10;
    addra = 32'd73408;
    dina = {96'd0, 16'd62625, 16'd15078, 16'd58413, 16'd46056, 16'd56936, 16'd51448, 16'd63794, 16'd20252, 16'd32985, 16'd15853}; // indx = 2294
    #10;
    addra = 32'd73440;
    dina = {96'd0, 16'd10334, 16'd39382, 16'd14482, 16'd49974, 16'd54553, 16'd30018, 16'd35134, 16'd28187, 16'd62668, 16'd63018}; // indx = 2295
    #10;
    addra = 32'd73472;
    dina = {96'd0, 16'd49327, 16'd6622, 16'd42613, 16'd7607, 16'd59485, 16'd28723, 16'd13444, 16'd59222, 16'd21481, 16'd9938}; // indx = 2296
    #10;
    addra = 32'd73504;
    dina = {96'd0, 16'd59822, 16'd927, 16'd18893, 16'd18348, 16'd65193, 16'd24977, 16'd16380, 16'd63294, 16'd3386, 16'd49839}; // indx = 2297
    #10;
    addra = 32'd73536;
    dina = {96'd0, 16'd27026, 16'd29633, 16'd46469, 16'd15297, 16'd47596, 16'd38199, 16'd18504, 16'd23245, 16'd14953, 16'd14349}; // indx = 2298
    #10;
    addra = 32'd73568;
    dina = {96'd0, 16'd36073, 16'd42620, 16'd35373, 16'd54192, 16'd54260, 16'd2024, 16'd40521, 16'd31256, 16'd38514, 16'd30989}; // indx = 2299
    #10;
    addra = 32'd73600;
    dina = {96'd0, 16'd56550, 16'd5688, 16'd53556, 16'd23610, 16'd2188, 16'd64457, 16'd5990, 16'd33142, 16'd26206, 16'd289}; // indx = 2300
    #10;
    addra = 32'd73632;
    dina = {96'd0, 16'd38625, 16'd18492, 16'd19698, 16'd16323, 16'd31360, 16'd18173, 16'd5309, 16'd13757, 16'd43640, 16'd26547}; // indx = 2301
    #10;
    addra = 32'd73664;
    dina = {96'd0, 16'd11778, 16'd19387, 16'd39562, 16'd47830, 16'd51766, 16'd5936, 16'd48144, 16'd18585, 16'd9840, 16'd43979}; // indx = 2302
    #10;
    addra = 32'd73696;
    dina = {96'd0, 16'd64465, 16'd15502, 16'd12086, 16'd32140, 16'd38069, 16'd10427, 16'd22675, 16'd12018, 16'd38301, 16'd16467}; // indx = 2303
    #10;
    addra = 32'd73728;
    dina = {96'd0, 16'd3235, 16'd11122, 16'd35268, 16'd265, 16'd43887, 16'd47156, 16'd45923, 16'd3806, 16'd60496, 16'd16729}; // indx = 2304
    #10;
    addra = 32'd73760;
    dina = {96'd0, 16'd53916, 16'd44403, 16'd45994, 16'd26193, 16'd41588, 16'd48986, 16'd63358, 16'd12025, 16'd42453, 16'd30340}; // indx = 2305
    #10;
    addra = 32'd73792;
    dina = {96'd0, 16'd8296, 16'd13501, 16'd58283, 16'd29842, 16'd15683, 16'd10834, 16'd2702, 16'd51557, 16'd13484, 16'd30770}; // indx = 2306
    #10;
    addra = 32'd73824;
    dina = {96'd0, 16'd49291, 16'd8790, 16'd1139, 16'd6639, 16'd50570, 16'd20132, 16'd59727, 16'd1919, 16'd51229, 16'd48007}; // indx = 2307
    #10;
    addra = 32'd73856;
    dina = {96'd0, 16'd14223, 16'd5385, 16'd10983, 16'd56784, 16'd26314, 16'd46747, 16'd36956, 16'd52866, 16'd46006, 16'd12298}; // indx = 2308
    #10;
    addra = 32'd73888;
    dina = {96'd0, 16'd30341, 16'd4973, 16'd6652, 16'd57716, 16'd41688, 16'd11254, 16'd6277, 16'd8160, 16'd63213, 16'd15908}; // indx = 2309
    #10;
    addra = 32'd73920;
    dina = {96'd0, 16'd64127, 16'd53331, 16'd30414, 16'd17219, 16'd28528, 16'd25555, 16'd21030, 16'd3643, 16'd27545, 16'd61362}; // indx = 2310
    #10;
    addra = 32'd73952;
    dina = {96'd0, 16'd52228, 16'd43947, 16'd33767, 16'd53858, 16'd55203, 16'd13380, 16'd37278, 16'd3968, 16'd31800, 16'd20438}; // indx = 2311
    #10;
    addra = 32'd73984;
    dina = {96'd0, 16'd13273, 16'd9597, 16'd407, 16'd20407, 16'd41153, 16'd61642, 16'd26251, 16'd36696, 16'd22738, 16'd44131}; // indx = 2312
    #10;
    addra = 32'd74016;
    dina = {96'd0, 16'd10768, 16'd41513, 16'd16888, 16'd29526, 16'd8520, 16'd64877, 16'd27024, 16'd28077, 16'd47432, 16'd3019}; // indx = 2313
    #10;
    addra = 32'd74048;
    dina = {96'd0, 16'd23078, 16'd57862, 16'd34360, 16'd36608, 16'd50217, 16'd26554, 16'd63404, 16'd17995, 16'd57336, 16'd50103}; // indx = 2314
    #10;
    addra = 32'd74080;
    dina = {96'd0, 16'd54251, 16'd29745, 16'd46505, 16'd28762, 16'd1944, 16'd5518, 16'd11667, 16'd64314, 16'd62918, 16'd10664}; // indx = 2315
    #10;
    addra = 32'd74112;
    dina = {96'd0, 16'd2716, 16'd59166, 16'd42494, 16'd9763, 16'd18571, 16'd8636, 16'd26834, 16'd4674, 16'd19484, 16'd10619}; // indx = 2316
    #10;
    addra = 32'd74144;
    dina = {96'd0, 16'd19914, 16'd65158, 16'd9031, 16'd19182, 16'd20865, 16'd51682, 16'd45598, 16'd61340, 16'd46783, 16'd59506}; // indx = 2317
    #10;
    addra = 32'd74176;
    dina = {96'd0, 16'd48585, 16'd17756, 16'd40886, 16'd56458, 16'd12278, 16'd6882, 16'd28056, 16'd47134, 16'd51699, 16'd35333}; // indx = 2318
    #10;
    addra = 32'd74208;
    dina = {96'd0, 16'd25344, 16'd13827, 16'd1421, 16'd57422, 16'd56689, 16'd2086, 16'd32881, 16'd52766, 16'd2664, 16'd785}; // indx = 2319
    #10;
    addra = 32'd74240;
    dina = {96'd0, 16'd21941, 16'd49830, 16'd55707, 16'd64310, 16'd33551, 16'd50360, 16'd55978, 16'd30171, 16'd22092, 16'd13506}; // indx = 2320
    #10;
    addra = 32'd74272;
    dina = {96'd0, 16'd20714, 16'd32636, 16'd37596, 16'd8054, 16'd5498, 16'd58160, 16'd42385, 16'd57687, 16'd42389, 16'd5169}; // indx = 2321
    #10;
    addra = 32'd74304;
    dina = {96'd0, 16'd31813, 16'd53416, 16'd30041, 16'd4912, 16'd51784, 16'd24865, 16'd38905, 16'd32359, 16'd54641, 16'd54532}; // indx = 2322
    #10;
    addra = 32'd74336;
    dina = {96'd0, 16'd52461, 16'd12590, 16'd26771, 16'd33162, 16'd53479, 16'd7705, 16'd30828, 16'd36972, 16'd26169, 16'd4434}; // indx = 2323
    #10;
    addra = 32'd74368;
    dina = {96'd0, 16'd56409, 16'd19802, 16'd54491, 16'd12933, 16'd64825, 16'd33865, 16'd5867, 16'd7968, 16'd49065, 16'd21209}; // indx = 2324
    #10;
    addra = 32'd74400;
    dina = {96'd0, 16'd64222, 16'd52097, 16'd6479, 16'd48807, 16'd20874, 16'd65420, 16'd8285, 16'd55721, 16'd43583, 16'd20353}; // indx = 2325
    #10;
    addra = 32'd74432;
    dina = {96'd0, 16'd5496, 16'd59556, 16'd37472, 16'd24296, 16'd57829, 16'd62738, 16'd3014, 16'd59912, 16'd20669, 16'd24249}; // indx = 2326
    #10;
    addra = 32'd74464;
    dina = {96'd0, 16'd16331, 16'd38694, 16'd3502, 16'd19050, 16'd36980, 16'd27465, 16'd54534, 16'd36295, 16'd18367, 16'd56789}; // indx = 2327
    #10;
    addra = 32'd74496;
    dina = {96'd0, 16'd23137, 16'd6197, 16'd11659, 16'd32317, 16'd40439, 16'd38355, 16'd37401, 16'd13585, 16'd59935, 16'd43451}; // indx = 2328
    #10;
    addra = 32'd74528;
    dina = {96'd0, 16'd121, 16'd39779, 16'd17178, 16'd32714, 16'd53147, 16'd40066, 16'd24111, 16'd45110, 16'd3778, 16'd52789}; // indx = 2329
    #10;
    addra = 32'd74560;
    dina = {96'd0, 16'd45361, 16'd4351, 16'd24889, 16'd24881, 16'd31049, 16'd1267, 16'd19827, 16'd23246, 16'd55485, 16'd63104}; // indx = 2330
    #10;
    addra = 32'd74592;
    dina = {96'd0, 16'd54414, 16'd23867, 16'd32995, 16'd31725, 16'd47258, 16'd22867, 16'd44218, 16'd27688, 16'd39031, 16'd2401}; // indx = 2331
    #10;
    addra = 32'd74624;
    dina = {96'd0, 16'd55154, 16'd60645, 16'd31808, 16'd35991, 16'd49563, 16'd4493, 16'd30208, 16'd64565, 16'd28720, 16'd1272}; // indx = 2332
    #10;
    addra = 32'd74656;
    dina = {96'd0, 16'd8348, 16'd32883, 16'd58944, 16'd38374, 16'd42137, 16'd23178, 16'd633, 16'd64426, 16'd19872, 16'd33804}; // indx = 2333
    #10;
    addra = 32'd74688;
    dina = {96'd0, 16'd12013, 16'd2138, 16'd9317, 16'd1362, 16'd46534, 16'd9212, 16'd16757, 16'd52320, 16'd15050, 16'd57058}; // indx = 2334
    #10;
    addra = 32'd74720;
    dina = {96'd0, 16'd40133, 16'd26286, 16'd38782, 16'd19659, 16'd29190, 16'd62902, 16'd2634, 16'd25685, 16'd8684, 16'd54503}; // indx = 2335
    #10;
    addra = 32'd74752;
    dina = {96'd0, 16'd51118, 16'd32139, 16'd57762, 16'd56215, 16'd37001, 16'd14410, 16'd47609, 16'd56763, 16'd4752, 16'd64983}; // indx = 2336
    #10;
    addra = 32'd74784;
    dina = {96'd0, 16'd25056, 16'd2633, 16'd15517, 16'd49367, 16'd23890, 16'd37203, 16'd50209, 16'd25078, 16'd58739, 16'd14782}; // indx = 2337
    #10;
    addra = 32'd74816;
    dina = {96'd0, 16'd8063, 16'd65148, 16'd63777, 16'd18649, 16'd39537, 16'd51742, 16'd8746, 16'd60191, 16'd37172, 16'd25517}; // indx = 2338
    #10;
    addra = 32'd74848;
    dina = {96'd0, 16'd19421, 16'd59073, 16'd44005, 16'd24436, 16'd28805, 16'd45562, 16'd27435, 16'd52513, 16'd26196, 16'd11562}; // indx = 2339
    #10;
    addra = 32'd74880;
    dina = {96'd0, 16'd27914, 16'd34999, 16'd52390, 16'd63870, 16'd54205, 16'd9099, 16'd2130, 16'd9093, 16'd50105, 16'd13885}; // indx = 2340
    #10;
    addra = 32'd74912;
    dina = {96'd0, 16'd23279, 16'd12370, 16'd54713, 16'd48930, 16'd25931, 16'd64135, 16'd15840, 16'd12886, 16'd63460, 16'd14082}; // indx = 2341
    #10;
    addra = 32'd74944;
    dina = {96'd0, 16'd57514, 16'd12402, 16'd44998, 16'd32507, 16'd8621, 16'd38393, 16'd55273, 16'd9322, 16'd40967, 16'd32711}; // indx = 2342
    #10;
    addra = 32'd74976;
    dina = {96'd0, 16'd60794, 16'd16183, 16'd34988, 16'd2002, 16'd20318, 16'd9104, 16'd48618, 16'd36998, 16'd57983, 16'd45416}; // indx = 2343
    #10;
    addra = 32'd75008;
    dina = {96'd0, 16'd60289, 16'd20715, 16'd32161, 16'd1386, 16'd34919, 16'd61487, 16'd41839, 16'd53983, 16'd15046, 16'd41196}; // indx = 2344
    #10;
    addra = 32'd75040;
    dina = {96'd0, 16'd35039, 16'd45783, 16'd19684, 16'd15635, 16'd45273, 16'd42413, 16'd51811, 16'd6421, 16'd34397, 16'd44704}; // indx = 2345
    #10;
    addra = 32'd75072;
    dina = {96'd0, 16'd2734, 16'd50966, 16'd20224, 16'd50462, 16'd47834, 16'd57845, 16'd60580, 16'd39873, 16'd10355, 16'd1889}; // indx = 2346
    #10;
    addra = 32'd75104;
    dina = {96'd0, 16'd58188, 16'd43702, 16'd26528, 16'd49771, 16'd48147, 16'd35532, 16'd5287, 16'd31883, 16'd51590, 16'd18672}; // indx = 2347
    #10;
    addra = 32'd75136;
    dina = {96'd0, 16'd5708, 16'd32459, 16'd7806, 16'd10989, 16'd42679, 16'd42121, 16'd61108, 16'd52766, 16'd60499, 16'd63595}; // indx = 2348
    #10;
    addra = 32'd75168;
    dina = {96'd0, 16'd43114, 16'd22162, 16'd27504, 16'd35626, 16'd3425, 16'd30078, 16'd7649, 16'd29693, 16'd607, 16'd16495}; // indx = 2349
    #10;
    addra = 32'd75200;
    dina = {96'd0, 16'd17444, 16'd37255, 16'd33504, 16'd43449, 16'd45312, 16'd39981, 16'd35173, 16'd14857, 16'd36288, 16'd37311}; // indx = 2350
    #10;
    addra = 32'd75232;
    dina = {96'd0, 16'd42891, 16'd55285, 16'd25095, 16'd27613, 16'd15026, 16'd52641, 16'd20400, 16'd1148, 16'd4980, 16'd34129}; // indx = 2351
    #10;
    addra = 32'd75264;
    dina = {96'd0, 16'd43957, 16'd62031, 16'd43141, 16'd62457, 16'd52575, 16'd23509, 16'd64819, 16'd31690, 16'd47283, 16'd46525}; // indx = 2352
    #10;
    addra = 32'd75296;
    dina = {96'd0, 16'd51678, 16'd36948, 16'd47537, 16'd44680, 16'd15622, 16'd33236, 16'd26724, 16'd58940, 16'd33377, 16'd5642}; // indx = 2353
    #10;
    addra = 32'd75328;
    dina = {96'd0, 16'd56118, 16'd19328, 16'd6386, 16'd50356, 16'd22881, 16'd35745, 16'd6602, 16'd36919, 16'd14630, 16'd42606}; // indx = 2354
    #10;
    addra = 32'd75360;
    dina = {96'd0, 16'd51267, 16'd12942, 16'd25960, 16'd3660, 16'd7512, 16'd37635, 16'd9809, 16'd1312, 16'd22790, 16'd54295}; // indx = 2355
    #10;
    addra = 32'd75392;
    dina = {96'd0, 16'd42434, 16'd33086, 16'd62742, 16'd5508, 16'd35587, 16'd49318, 16'd18778, 16'd52429, 16'd15621, 16'd55957}; // indx = 2356
    #10;
    addra = 32'd75424;
    dina = {96'd0, 16'd15414, 16'd25668, 16'd64274, 16'd1823, 16'd53777, 16'd21749, 16'd64204, 16'd38719, 16'd55415, 16'd57236}; // indx = 2357
    #10;
    addra = 32'd75456;
    dina = {96'd0, 16'd12832, 16'd45351, 16'd35747, 16'd46929, 16'd42762, 16'd1535, 16'd15145, 16'd54756, 16'd22736, 16'd43783}; // indx = 2358
    #10;
    addra = 32'd75488;
    dina = {96'd0, 16'd63736, 16'd48480, 16'd42854, 16'd35869, 16'd17140, 16'd21057, 16'd50490, 16'd15822, 16'd65100, 16'd29253}; // indx = 2359
    #10;
    addra = 32'd75520;
    dina = {96'd0, 16'd26400, 16'd51113, 16'd55745, 16'd470, 16'd46656, 16'd62243, 16'd9912, 16'd1412, 16'd40232, 16'd373}; // indx = 2360
    #10;
    addra = 32'd75552;
    dina = {96'd0, 16'd45394, 16'd25743, 16'd10064, 16'd31229, 16'd31300, 16'd42740, 16'd26709, 16'd60598, 16'd36962, 16'd35413}; // indx = 2361
    #10;
    addra = 32'd75584;
    dina = {96'd0, 16'd53550, 16'd45505, 16'd11764, 16'd46497, 16'd20494, 16'd40171, 16'd10177, 16'd65246, 16'd56446, 16'd41214}; // indx = 2362
    #10;
    addra = 32'd75616;
    dina = {96'd0, 16'd25141, 16'd64205, 16'd52494, 16'd28772, 16'd61805, 16'd23537, 16'd13739, 16'd8661, 16'd37312, 16'd64}; // indx = 2363
    #10;
    addra = 32'd75648;
    dina = {96'd0, 16'd57325, 16'd59575, 16'd58745, 16'd17846, 16'd49895, 16'd38624, 16'd2876, 16'd44427, 16'd6404, 16'd52269}; // indx = 2364
    #10;
    addra = 32'd75680;
    dina = {96'd0, 16'd36173, 16'd63042, 16'd32127, 16'd16049, 16'd47199, 16'd32152, 16'd49925, 16'd3550, 16'd26757, 16'd1953}; // indx = 2365
    #10;
    addra = 32'd75712;
    dina = {96'd0, 16'd5355, 16'd17014, 16'd59488, 16'd18710, 16'd27657, 16'd30506, 16'd17914, 16'd54681, 16'd45714, 16'd61452}; // indx = 2366
    #10;
    addra = 32'd75744;
    dina = {96'd0, 16'd19098, 16'd59806, 16'd24406, 16'd35228, 16'd2627, 16'd34802, 16'd53602, 16'd48144, 16'd7400, 16'd38662}; // indx = 2367
    #10;
    addra = 32'd75776;
    dina = {96'd0, 16'd64066, 16'd12332, 16'd20431, 16'd26514, 16'd57137, 16'd60293, 16'd63518, 16'd547, 16'd30985, 16'd31686}; // indx = 2368
    #10;
    addra = 32'd75808;
    dina = {96'd0, 16'd5864, 16'd54966, 16'd63300, 16'd2577, 16'd8420, 16'd46411, 16'd58270, 16'd53424, 16'd46647, 16'd30178}; // indx = 2369
    #10;
    addra = 32'd75840;
    dina = {96'd0, 16'd21077, 16'd7716, 16'd34127, 16'd62959, 16'd37970, 16'd35236, 16'd10373, 16'd51022, 16'd41573, 16'd7699}; // indx = 2370
    #10;
    addra = 32'd75872;
    dina = {96'd0, 16'd35125, 16'd10213, 16'd2147, 16'd37736, 16'd19445, 16'd46425, 16'd15405, 16'd4025, 16'd64917, 16'd38912}; // indx = 2371
    #10;
    addra = 32'd75904;
    dina = {96'd0, 16'd21514, 16'd40775, 16'd33877, 16'd28359, 16'd34121, 16'd7163, 16'd8631, 16'd46348, 16'd48689, 16'd51435}; // indx = 2372
    #10;
    addra = 32'd75936;
    dina = {96'd0, 16'd52858, 16'd22303, 16'd9316, 16'd11273, 16'd38525, 16'd4746, 16'd40976, 16'd48446, 16'd53184, 16'd3749}; // indx = 2373
    #10;
    addra = 32'd75968;
    dina = {96'd0, 16'd49861, 16'd63129, 16'd23809, 16'd545, 16'd12722, 16'd41114, 16'd23782, 16'd21787, 16'd56635, 16'd49974}; // indx = 2374
    #10;
    addra = 32'd76000;
    dina = {96'd0, 16'd4315, 16'd38483, 16'd19890, 16'd15676, 16'd34331, 16'd7123, 16'd4082, 16'd55590, 16'd42728, 16'd61898}; // indx = 2375
    #10;
    addra = 32'd76032;
    dina = {96'd0, 16'd52846, 16'd20338, 16'd41340, 16'd9485, 16'd40828, 16'd25245, 16'd17826, 16'd60984, 16'd37154, 16'd35888}; // indx = 2376
    #10;
    addra = 32'd76064;
    dina = {96'd0, 16'd49841, 16'd26652, 16'd56699, 16'd10450, 16'd62486, 16'd33089, 16'd42330, 16'd35642, 16'd2844, 16'd17904}; // indx = 2377
    #10;
    addra = 32'd76096;
    dina = {96'd0, 16'd22435, 16'd50662, 16'd15232, 16'd38260, 16'd26714, 16'd6490, 16'd59641, 16'd11329, 16'd31069, 16'd11077}; // indx = 2378
    #10;
    addra = 32'd76128;
    dina = {96'd0, 16'd56648, 16'd48218, 16'd12221, 16'd49834, 16'd12623, 16'd24044, 16'd42616, 16'd4934, 16'd39150, 16'd27102}; // indx = 2379
    #10;
    addra = 32'd76160;
    dina = {96'd0, 16'd55548, 16'd28577, 16'd29358, 16'd51590, 16'd23205, 16'd31102, 16'd32002, 16'd25728, 16'd4833, 16'd63919}; // indx = 2380
    #10;
    addra = 32'd76192;
    dina = {96'd0, 16'd50401, 16'd19084, 16'd32345, 16'd9521, 16'd8146, 16'd34565, 16'd5633, 16'd32448, 16'd60501, 16'd33907}; // indx = 2381
    #10;
    addra = 32'd76224;
    dina = {96'd0, 16'd19920, 16'd44250, 16'd9127, 16'd45121, 16'd14142, 16'd16106, 16'd51101, 16'd1806, 16'd18330, 16'd54575}; // indx = 2382
    #10;
    addra = 32'd76256;
    dina = {96'd0, 16'd21084, 16'd14274, 16'd18052, 16'd41398, 16'd26906, 16'd42220, 16'd37846, 16'd22481, 16'd39794, 16'd21583}; // indx = 2383
    #10;
    addra = 32'd76288;
    dina = {96'd0, 16'd44411, 16'd47801, 16'd39931, 16'd28147, 16'd62074, 16'd43637, 16'd23084, 16'd57915, 16'd19116, 16'd52489}; // indx = 2384
    #10;
    addra = 32'd76320;
    dina = {96'd0, 16'd35660, 16'd40011, 16'd5034, 16'd57952, 16'd44378, 16'd18848, 16'd27162, 16'd48789, 16'd38518, 16'd59112}; // indx = 2385
    #10;
    addra = 32'd76352;
    dina = {96'd0, 16'd31567, 16'd34150, 16'd7045, 16'd56222, 16'd29572, 16'd31618, 16'd65313, 16'd38001, 16'd16262, 16'd10137}; // indx = 2386
    #10;
    addra = 32'd76384;
    dina = {96'd0, 16'd64116, 16'd16195, 16'd36415, 16'd27475, 16'd32822, 16'd44785, 16'd50312, 16'd4702, 16'd31610, 16'd55703}; // indx = 2387
    #10;
    addra = 32'd76416;
    dina = {96'd0, 16'd13573, 16'd27839, 16'd8831, 16'd51778, 16'd47392, 16'd48770, 16'd30886, 16'd14582, 16'd49218, 16'd55388}; // indx = 2388
    #10;
    addra = 32'd76448;
    dina = {96'd0, 16'd43537, 16'd34911, 16'd12402, 16'd9530, 16'd30829, 16'd48482, 16'd36280, 16'd16903, 16'd19236, 16'd11776}; // indx = 2389
    #10;
    addra = 32'd76480;
    dina = {96'd0, 16'd57657, 16'd11452, 16'd64974, 16'd12615, 16'd64234, 16'd25735, 16'd57819, 16'd8908, 16'd54601, 16'd1701}; // indx = 2390
    #10;
    addra = 32'd76512;
    dina = {96'd0, 16'd23344, 16'd25645, 16'd915, 16'd48900, 16'd27419, 16'd2645, 16'd48986, 16'd10322, 16'd16695, 16'd55058}; // indx = 2391
    #10;
    addra = 32'd76544;
    dina = {96'd0, 16'd29171, 16'd30293, 16'd15876, 16'd297, 16'd25512, 16'd11060, 16'd50381, 16'd53548, 16'd59943, 16'd22140}; // indx = 2392
    #10;
    addra = 32'd76576;
    dina = {96'd0, 16'd44262, 16'd42982, 16'd40835, 16'd12206, 16'd4196, 16'd2578, 16'd15554, 16'd41504, 16'd29873, 16'd53931}; // indx = 2393
    #10;
    addra = 32'd76608;
    dina = {96'd0, 16'd23109, 16'd50547, 16'd55412, 16'd21677, 16'd33519, 16'd28139, 16'd52830, 16'd18539, 16'd46969, 16'd22496}; // indx = 2394
    #10;
    addra = 32'd76640;
    dina = {96'd0, 16'd48225, 16'd6912, 16'd57133, 16'd47608, 16'd55249, 16'd19994, 16'd46272, 16'd55109, 16'd56397, 16'd19883}; // indx = 2395
    #10;
    addra = 32'd76672;
    dina = {96'd0, 16'd34754, 16'd44358, 16'd32009, 16'd33384, 16'd8939, 16'd8252, 16'd64644, 16'd43688, 16'd43877, 16'd46392}; // indx = 2396
    #10;
    addra = 32'd76704;
    dina = {96'd0, 16'd9045, 16'd19252, 16'd23263, 16'd11602, 16'd58524, 16'd58325, 16'd44667, 16'd63106, 16'd20687, 16'd58210}; // indx = 2397
    #10;
    addra = 32'd76736;
    dina = {96'd0, 16'd44737, 16'd11855, 16'd41112, 16'd44288, 16'd52087, 16'd20697, 16'd63534, 16'd29423, 16'd46662, 16'd44795}; // indx = 2398
    #10;
    addra = 32'd76768;
    dina = {96'd0, 16'd33913, 16'd41900, 16'd62929, 16'd12156, 16'd44554, 16'd7116, 16'd57178, 16'd6466, 16'd401, 16'd7311}; // indx = 2399
    #10;
    addra = 32'd76800;
    dina = {96'd0, 16'd48928, 16'd43763, 16'd33806, 16'd62046, 16'd9074, 16'd2885, 16'd51492, 16'd24828, 16'd39024, 16'd36616}; // indx = 2400
    #10;
    addra = 32'd76832;
    dina = {96'd0, 16'd21906, 16'd11295, 16'd21643, 16'd10636, 16'd60748, 16'd7061, 16'd50389, 16'd14200, 16'd42395, 16'd26264}; // indx = 2401
    #10;
    addra = 32'd76864;
    dina = {96'd0, 16'd21442, 16'd21418, 16'd4939, 16'd62918, 16'd31845, 16'd45170, 16'd33223, 16'd13901, 16'd5918, 16'd39764}; // indx = 2402
    #10;
    addra = 32'd76896;
    dina = {96'd0, 16'd11384, 16'd3125, 16'd12065, 16'd58130, 16'd46455, 16'd13747, 16'd26514, 16'd32505, 16'd49673, 16'd18429}; // indx = 2403
    #10;
    addra = 32'd76928;
    dina = {96'd0, 16'd15495, 16'd43049, 16'd57949, 16'd16064, 16'd45210, 16'd16414, 16'd20676, 16'd49481, 16'd62834, 16'd36806}; // indx = 2404
    #10;
    addra = 32'd76960;
    dina = {96'd0, 16'd58330, 16'd43552, 16'd43353, 16'd8520, 16'd14873, 16'd56411, 16'd5408, 16'd3148, 16'd64212, 16'd6352}; // indx = 2405
    #10;
    addra = 32'd76992;
    dina = {96'd0, 16'd57682, 16'd3236, 16'd61136, 16'd44327, 16'd5890, 16'd43680, 16'd50367, 16'd13831, 16'd18970, 16'd47647}; // indx = 2406
    #10;
    addra = 32'd77024;
    dina = {96'd0, 16'd55475, 16'd37479, 16'd60493, 16'd11065, 16'd20128, 16'd15312, 16'd16317, 16'd65059, 16'd25803, 16'd61269}; // indx = 2407
    #10;
    addra = 32'd77056;
    dina = {96'd0, 16'd39832, 16'd47211, 16'd26632, 16'd9878, 16'd52755, 16'd47330, 16'd8120, 16'd3718, 16'd3936, 16'd7249}; // indx = 2408
    #10;
    addra = 32'd77088;
    dina = {96'd0, 16'd34765, 16'd49785, 16'd22266, 16'd20744, 16'd41625, 16'd46092, 16'd38777, 16'd38192, 16'd11197, 16'd15391}; // indx = 2409
    #10;
    addra = 32'd77120;
    dina = {96'd0, 16'd21293, 16'd23494, 16'd5804, 16'd54675, 16'd56335, 16'd16698, 16'd11583, 16'd43389, 16'd45455, 16'd57988}; // indx = 2410
    #10;
    addra = 32'd77152;
    dina = {96'd0, 16'd34298, 16'd53091, 16'd3701, 16'd2807, 16'd13059, 16'd55686, 16'd27493, 16'd6428, 16'd13191, 16'd56760}; // indx = 2411
    #10;
    addra = 32'd77184;
    dina = {96'd0, 16'd63857, 16'd17951, 16'd8544, 16'd64488, 16'd64802, 16'd59343, 16'd55498, 16'd7841, 16'd33498, 16'd20724}; // indx = 2412
    #10;
    addra = 32'd77216;
    dina = {96'd0, 16'd62571, 16'd38259, 16'd13731, 16'd47768, 16'd33016, 16'd8700, 16'd895, 16'd47525, 16'd13853, 16'd4197}; // indx = 2413
    #10;
    addra = 32'd77248;
    dina = {96'd0, 16'd40770, 16'd63768, 16'd57033, 16'd46113, 16'd29605, 16'd19543, 16'd48710, 16'd31264, 16'd32814, 16'd25399}; // indx = 2414
    #10;
    addra = 32'd77280;
    dina = {96'd0, 16'd29193, 16'd56024, 16'd31898, 16'd3855, 16'd30963, 16'd26944, 16'd34615, 16'd20354, 16'd8042, 16'd55000}; // indx = 2415
    #10;
    addra = 32'd77312;
    dina = {96'd0, 16'd32879, 16'd26278, 16'd50557, 16'd35131, 16'd33619, 16'd16348, 16'd37057, 16'd54127, 16'd23790, 16'd35812}; // indx = 2416
    #10;
    addra = 32'd77344;
    dina = {96'd0, 16'd36183, 16'd63195, 16'd19292, 16'd33278, 16'd49749, 16'd59829, 16'd4217, 16'd32013, 16'd883, 16'd9002}; // indx = 2417
    #10;
    addra = 32'd77376;
    dina = {96'd0, 16'd57279, 16'd12221, 16'd51947, 16'd60563, 16'd24453, 16'd36958, 16'd17542, 16'd60369, 16'd56666, 16'd37967}; // indx = 2418
    #10;
    addra = 32'd77408;
    dina = {96'd0, 16'd33807, 16'd37178, 16'd27018, 16'd12614, 16'd354, 16'd32757, 16'd50107, 16'd18262, 16'd712, 16'd45892}; // indx = 2419
    #10;
    addra = 32'd77440;
    dina = {96'd0, 16'd40980, 16'd31761, 16'd19979, 16'd26103, 16'd28164, 16'd16057, 16'd4711, 16'd34299, 16'd29823, 16'd31883}; // indx = 2420
    #10;
    addra = 32'd77472;
    dina = {96'd0, 16'd10730, 16'd37794, 16'd39555, 16'd41830, 16'd47194, 16'd62017, 16'd18635, 16'd41103, 16'd42055, 16'd51362}; // indx = 2421
    #10;
    addra = 32'd77504;
    dina = {96'd0, 16'd50637, 16'd14251, 16'd44381, 16'd45909, 16'd22681, 16'd17422, 16'd49231, 16'd10273, 16'd51334, 16'd54604}; // indx = 2422
    #10;
    addra = 32'd77536;
    dina = {96'd0, 16'd44060, 16'd44061, 16'd48188, 16'd30418, 16'd45147, 16'd3846, 16'd54988, 16'd9534, 16'd29909, 16'd45057}; // indx = 2423
    #10;
    addra = 32'd77568;
    dina = {96'd0, 16'd62366, 16'd13403, 16'd14013, 16'd27830, 16'd35733, 16'd15227, 16'd25956, 16'd58259, 16'd54058, 16'd43557}; // indx = 2424
    #10;
    addra = 32'd77600;
    dina = {96'd0, 16'd54020, 16'd31651, 16'd15305, 16'd36683, 16'd31723, 16'd57583, 16'd4249, 16'd47139, 16'd40810, 16'd64808}; // indx = 2425
    #10;
    addra = 32'd77632;
    dina = {96'd0, 16'd9348, 16'd40821, 16'd28077, 16'd18540, 16'd31157, 16'd14164, 16'd10054, 16'd56264, 16'd37113, 16'd65025}; // indx = 2426
    #10;
    addra = 32'd77664;
    dina = {96'd0, 16'd45628, 16'd22185, 16'd40765, 16'd36819, 16'd8748, 16'd54936, 16'd43119, 16'd10203, 16'd19451, 16'd32471}; // indx = 2427
    #10;
    addra = 32'd77696;
    dina = {96'd0, 16'd3038, 16'd57438, 16'd45434, 16'd37011, 16'd26271, 16'd28440, 16'd5535, 16'd1677, 16'd63509, 16'd4532}; // indx = 2428
    #10;
    addra = 32'd77728;
    dina = {96'd0, 16'd26282, 16'd55720, 16'd37409, 16'd6507, 16'd6599, 16'd43634, 16'd33387, 16'd3254, 16'd58743, 16'd43797}; // indx = 2429
    #10;
    addra = 32'd77760;
    dina = {96'd0, 16'd5416, 16'd41879, 16'd44299, 16'd13282, 16'd23453, 16'd40509, 16'd46271, 16'd49888, 16'd41459, 16'd48981}; // indx = 2430
    #10;
    addra = 32'd77792;
    dina = {96'd0, 16'd17584, 16'd32401, 16'd40523, 16'd15141, 16'd39386, 16'd3243, 16'd24993, 16'd24341, 16'd4593, 16'd19413}; // indx = 2431
    #10;
    addra = 32'd77824;
    dina = {96'd0, 16'd44800, 16'd60338, 16'd63394, 16'd59112, 16'd55748, 16'd4773, 16'd25471, 16'd29314, 16'd37040, 16'd44306}; // indx = 2432
    #10;
    addra = 32'd77856;
    dina = {96'd0, 16'd31420, 16'd61231, 16'd57138, 16'd7878, 16'd640, 16'd47294, 16'd35606, 16'd17862, 16'd33322, 16'd63615}; // indx = 2433
    #10;
    addra = 32'd77888;
    dina = {96'd0, 16'd44350, 16'd63262, 16'd48532, 16'd55803, 16'd13282, 16'd58770, 16'd5284, 16'd16365, 16'd8629, 16'd42241}; // indx = 2434
    #10;
    addra = 32'd77920;
    dina = {96'd0, 16'd15741, 16'd62981, 16'd19324, 16'd45074, 16'd49891, 16'd61624, 16'd29867, 16'd23011, 16'd41093, 16'd31164}; // indx = 2435
    #10;
    addra = 32'd77952;
    dina = {96'd0, 16'd36508, 16'd17980, 16'd4062, 16'd4148, 16'd4226, 16'd32533, 16'd47564, 16'd31209, 16'd56914, 16'd5058}; // indx = 2436
    #10;
    addra = 32'd77984;
    dina = {96'd0, 16'd63670, 16'd61207, 16'd64090, 16'd63891, 16'd47722, 16'd33627, 16'd5310, 16'd57214, 16'd2674, 16'd27883}; // indx = 2437
    #10;
    addra = 32'd78016;
    dina = {96'd0, 16'd39731, 16'd39944, 16'd29132, 16'd43436, 16'd39885, 16'd24512, 16'd62842, 16'd46631, 16'd57558, 16'd45846}; // indx = 2438
    #10;
    addra = 32'd78048;
    dina = {96'd0, 16'd24034, 16'd30515, 16'd19028, 16'd14455, 16'd18647, 16'd14006, 16'd9310, 16'd51455, 16'd29477, 16'd25422}; // indx = 2439
    #10;
    addra = 32'd78080;
    dina = {96'd0, 16'd43227, 16'd40486, 16'd7345, 16'd29687, 16'd47216, 16'd20468, 16'd10749, 16'd31380, 16'd65227, 16'd19798}; // indx = 2440
    #10;
    addra = 32'd78112;
    dina = {96'd0, 16'd53398, 16'd32162, 16'd3780, 16'd38628, 16'd44582, 16'd33613, 16'd29200, 16'd59737, 16'd58798, 16'd23380}; // indx = 2441
    #10;
    addra = 32'd78144;
    dina = {96'd0, 16'd22996, 16'd41008, 16'd46885, 16'd21766, 16'd1210, 16'd50880, 16'd27602, 16'd38243, 16'd31726, 16'd45624}; // indx = 2442
    #10;
    addra = 32'd78176;
    dina = {96'd0, 16'd8664, 16'd38662, 16'd9482, 16'd7627, 16'd30873, 16'd3787, 16'd31557, 16'd23214, 16'd27373, 16'd63412}; // indx = 2443
    #10;
    addra = 32'd78208;
    dina = {96'd0, 16'd61180, 16'd8760, 16'd15349, 16'd51411, 16'd61806, 16'd17014, 16'd50176, 16'd35702, 16'd30364, 16'd44674}; // indx = 2444
    #10;
    addra = 32'd78240;
    dina = {96'd0, 16'd18487, 16'd652, 16'd2683, 16'd9294, 16'd57454, 16'd30673, 16'd49010, 16'd59606, 16'd42453, 16'd29379}; // indx = 2445
    #10;
    addra = 32'd78272;
    dina = {96'd0, 16'd54057, 16'd42515, 16'd5789, 16'd38881, 16'd45096, 16'd50590, 16'd18671, 16'd52801, 16'd34167, 16'd37631}; // indx = 2446
    #10;
    addra = 32'd78304;
    dina = {96'd0, 16'd44892, 16'd1674, 16'd40532, 16'd32676, 16'd47634, 16'd16345, 16'd43823, 16'd41752, 16'd40120, 16'd36469}; // indx = 2447
    #10;
    addra = 32'd78336;
    dina = {96'd0, 16'd11017, 16'd58905, 16'd18139, 16'd50394, 16'd3638, 16'd20051, 16'd5727, 16'd31237, 16'd32312, 16'd56426}; // indx = 2448
    #10;
    addra = 32'd78368;
    dina = {96'd0, 16'd21126, 16'd20871, 16'd45043, 16'd48524, 16'd30229, 16'd64768, 16'd54383, 16'd6496, 16'd8367, 16'd54539}; // indx = 2449
    #10;
    addra = 32'd78400;
    dina = {96'd0, 16'd61283, 16'd46174, 16'd25890, 16'd42665, 16'd5670, 16'd51935, 16'd26704, 16'd13748, 16'd39135, 16'd27409}; // indx = 2450
    #10;
    addra = 32'd78432;
    dina = {96'd0, 16'd12594, 16'd8628, 16'd39872, 16'd51495, 16'd21579, 16'd51346, 16'd24786, 16'd31076, 16'd13321, 16'd31850}; // indx = 2451
    #10;
    addra = 32'd78464;
    dina = {96'd0, 16'd4896, 16'd52192, 16'd16320, 16'd45770, 16'd41096, 16'd45205, 16'd25093, 16'd12980, 16'd45473, 16'd48646}; // indx = 2452
    #10;
    addra = 32'd78496;
    dina = {96'd0, 16'd34792, 16'd944, 16'd46424, 16'd15856, 16'd61912, 16'd59185, 16'd50546, 16'd48970, 16'd5422, 16'd22884}; // indx = 2453
    #10;
    addra = 32'd78528;
    dina = {96'd0, 16'd2919, 16'd26376, 16'd61592, 16'd48900, 16'd30394, 16'd17536, 16'd63846, 16'd61497, 16'd10613, 16'd43689}; // indx = 2454
    #10;
    addra = 32'd78560;
    dina = {96'd0, 16'd51378, 16'd28082, 16'd30395, 16'd35992, 16'd46865, 16'd12893, 16'd31653, 16'd29100, 16'd59034, 16'd22015}; // indx = 2455
    #10;
    addra = 32'd78592;
    dina = {96'd0, 16'd40064, 16'd14633, 16'd47128, 16'd32012, 16'd58668, 16'd60413, 16'd53499, 16'd61274, 16'd26059, 16'd25993}; // indx = 2456
    #10;
    addra = 32'd78624;
    dina = {96'd0, 16'd3363, 16'd397, 16'd30001, 16'd64362, 16'd22063, 16'd58851, 16'd59592, 16'd47118, 16'd38259, 16'd9552}; // indx = 2457
    #10;
    addra = 32'd78656;
    dina = {96'd0, 16'd25583, 16'd33414, 16'd9397, 16'd62960, 16'd21411, 16'd19803, 16'd45681, 16'd1203, 16'd24744, 16'd2221}; // indx = 2458
    #10;
    addra = 32'd78688;
    dina = {96'd0, 16'd8847, 16'd54259, 16'd9633, 16'd35912, 16'd11266, 16'd49318, 16'd55586, 16'd13926, 16'd47601, 16'd37243}; // indx = 2459
    #10;
    addra = 32'd78720;
    dina = {96'd0, 16'd63978, 16'd7043, 16'd38153, 16'd53767, 16'd18438, 16'd45928, 16'd3402, 16'd42460, 16'd7871, 16'd57227}; // indx = 2460
    #10;
    addra = 32'd78752;
    dina = {96'd0, 16'd9410, 16'd33993, 16'd8054, 16'd14956, 16'd25225, 16'd1600, 16'd61098, 16'd1721, 16'd31890, 16'd27897}; // indx = 2461
    #10;
    addra = 32'd78784;
    dina = {96'd0, 16'd54963, 16'd14451, 16'd40666, 16'd52233, 16'd19822, 16'd26159, 16'd21708, 16'd4053, 16'd27109, 16'd29206}; // indx = 2462
    #10;
    addra = 32'd78816;
    dina = {96'd0, 16'd51430, 16'd34727, 16'd50777, 16'd20593, 16'd49004, 16'd17891, 16'd29236, 16'd42083, 16'd54043, 16'd6077}; // indx = 2463
    #10;
    addra = 32'd78848;
    dina = {96'd0, 16'd60829, 16'd34988, 16'd30166, 16'd28010, 16'd18962, 16'd60411, 16'd48188, 16'd668, 16'd60524, 16'd57931}; // indx = 2464
    #10;
    addra = 32'd78880;
    dina = {96'd0, 16'd64201, 16'd9395, 16'd19907, 16'd51932, 16'd42866, 16'd14376, 16'd45281, 16'd60500, 16'd55643, 16'd21390}; // indx = 2465
    #10;
    addra = 32'd78912;
    dina = {96'd0, 16'd30372, 16'd37418, 16'd47201, 16'd63848, 16'd9103, 16'd60274, 16'd3689, 16'd25462, 16'd32983, 16'd41774}; // indx = 2466
    #10;
    addra = 32'd78944;
    dina = {96'd0, 16'd53634, 16'd13669, 16'd38156, 16'd41662, 16'd56026, 16'd18553, 16'd58761, 16'd35392, 16'd54939, 16'd37182}; // indx = 2467
    #10;
    addra = 32'd78976;
    dina = {96'd0, 16'd37471, 16'd74, 16'd25470, 16'd21615, 16'd31957, 16'd20951, 16'd12252, 16'd3477, 16'd20097, 16'd41464}; // indx = 2468
    #10;
    addra = 32'd79008;
    dina = {96'd0, 16'd3952, 16'd52694, 16'd6422, 16'd4845, 16'd39004, 16'd10345, 16'd27561, 16'd6574, 16'd39850, 16'd49085}; // indx = 2469
    #10;
    addra = 32'd79040;
    dina = {96'd0, 16'd61264, 16'd49662, 16'd37740, 16'd13478, 16'd40059, 16'd40346, 16'd25689, 16'd29148, 16'd19198, 16'd2222}; // indx = 2470
    #10;
    addra = 32'd79072;
    dina = {96'd0, 16'd9686, 16'd8174, 16'd7807, 16'd22533, 16'd47710, 16'd30564, 16'd18403, 16'd41025, 16'd49341, 16'd34407}; // indx = 2471
    #10;
    addra = 32'd79104;
    dina = {96'd0, 16'd63814, 16'd5472, 16'd16212, 16'd63342, 16'd19543, 16'd27382, 16'd2513, 16'd59158, 16'd24352, 16'd10173}; // indx = 2472
    #10;
    addra = 32'd79136;
    dina = {96'd0, 16'd19393, 16'd32086, 16'd64470, 16'd49164, 16'd34181, 16'd12069, 16'd4214, 16'd36891, 16'd42760, 16'd57451}; // indx = 2473
    #10;
    addra = 32'd79168;
    dina = {96'd0, 16'd41, 16'd40791, 16'd56893, 16'd7420, 16'd34206, 16'd50052, 16'd46332, 16'd50110, 16'd36902, 16'd53555}; // indx = 2474
    #10;
    addra = 32'd79200;
    dina = {96'd0, 16'd28443, 16'd51166, 16'd33264, 16'd46779, 16'd44151, 16'd51052, 16'd13271, 16'd39504, 16'd6464, 16'd40118}; // indx = 2475
    #10;
    addra = 32'd79232;
    dina = {96'd0, 16'd9587, 16'd36090, 16'd64996, 16'd8958, 16'd4732, 16'd57169, 16'd13996, 16'd48124, 16'd44126, 16'd53831}; // indx = 2476
    #10;
    addra = 32'd79264;
    dina = {96'd0, 16'd48614, 16'd32514, 16'd44752, 16'd4463, 16'd8481, 16'd63344, 16'd49718, 16'd15446, 16'd41781, 16'd25030}; // indx = 2477
    #10;
    addra = 32'd79296;
    dina = {96'd0, 16'd8105, 16'd4524, 16'd9725, 16'd26438, 16'd13311, 16'd62293, 16'd226, 16'd55081, 16'd23017, 16'd22483}; // indx = 2478
    #10;
    addra = 32'd79328;
    dina = {96'd0, 16'd55273, 16'd20452, 16'd12246, 16'd21644, 16'd27122, 16'd53076, 16'd7537, 16'd31500, 16'd17822, 16'd57831}; // indx = 2479
    #10;
    addra = 32'd79360;
    dina = {96'd0, 16'd26096, 16'd37305, 16'd31282, 16'd65239, 16'd17650, 16'd40695, 16'd22142, 16'd62230, 16'd48556, 16'd34922}; // indx = 2480
    #10;
    addra = 32'd79392;
    dina = {96'd0, 16'd27577, 16'd3233, 16'd16260, 16'd32542, 16'd61597, 16'd18799, 16'd10088, 16'd28200, 16'd40095, 16'd62279}; // indx = 2481
    #10;
    addra = 32'd79424;
    dina = {96'd0, 16'd37374, 16'd4702, 16'd28485, 16'd1712, 16'd59279, 16'd14415, 16'd26061, 16'd12665, 16'd27228, 16'd6492}; // indx = 2482
    #10;
    addra = 32'd79456;
    dina = {96'd0, 16'd34427, 16'd58768, 16'd33300, 16'd18286, 16'd54934, 16'd41608, 16'd42724, 16'd52408, 16'd63792, 16'd9830}; // indx = 2483
    #10;
    addra = 32'd79488;
    dina = {96'd0, 16'd55361, 16'd37211, 16'd51655, 16'd35603, 16'd14947, 16'd44664, 16'd48361, 16'd7946, 16'd51837, 16'd42908}; // indx = 2484
    #10;
    addra = 32'd79520;
    dina = {96'd0, 16'd6664, 16'd45970, 16'd16007, 16'd61923, 16'd12227, 16'd43982, 16'd62825, 16'd27905, 16'd34399, 16'd64565}; // indx = 2485
    #10;
    addra = 32'd79552;
    dina = {96'd0, 16'd59013, 16'd3630, 16'd64675, 16'd22342, 16'd14437, 16'd5348, 16'd57370, 16'd15085, 16'd52905, 16'd41613}; // indx = 2486
    #10;
    addra = 32'd79584;
    dina = {96'd0, 16'd59267, 16'd61605, 16'd29974, 16'd6057, 16'd18595, 16'd44203, 16'd60156, 16'd49151, 16'd29172, 16'd56756}; // indx = 2487
    #10;
    addra = 32'd79616;
    dina = {96'd0, 16'd21481, 16'd34723, 16'd14602, 16'd65506, 16'd12174, 16'd24317, 16'd6130, 16'd33132, 16'd54213, 16'd35135}; // indx = 2488
    #10;
    addra = 32'd79648;
    dina = {96'd0, 16'd22696, 16'd41983, 16'd65176, 16'd15748, 16'd32077, 16'd53198, 16'd44175, 16'd61004, 16'd63832, 16'd39457}; // indx = 2489
    #10;
    addra = 32'd79680;
    dina = {96'd0, 16'd63433, 16'd57083, 16'd43879, 16'd44644, 16'd12244, 16'd15908, 16'd12447, 16'd10793, 16'd2029, 16'd18795}; // indx = 2490
    #10;
    addra = 32'd79712;
    dina = {96'd0, 16'd26072, 16'd52960, 16'd48335, 16'd24161, 16'd28282, 16'd58590, 16'd60775, 16'd29857, 16'd15960, 16'd32574}; // indx = 2491
    #10;
    addra = 32'd79744;
    dina = {96'd0, 16'd49458, 16'd15565, 16'd59026, 16'd11766, 16'd46116, 16'd45011, 16'd27434, 16'd33644, 16'd34081, 16'd60184}; // indx = 2492
    #10;
    addra = 32'd79776;
    dina = {96'd0, 16'd64871, 16'd37232, 16'd65467, 16'd37431, 16'd62095, 16'd55148, 16'd10372, 16'd56466, 16'd58603, 16'd64437}; // indx = 2493
    #10;
    addra = 32'd79808;
    dina = {96'd0, 16'd63611, 16'd35952, 16'd30095, 16'd57706, 16'd62659, 16'd50302, 16'd45567, 16'd34607, 16'd11379, 16'd3750}; // indx = 2494
    #10;
    addra = 32'd79840;
    dina = {96'd0, 16'd664, 16'd47048, 16'd22495, 16'd63012, 16'd51874, 16'd58980, 16'd51525, 16'd40982, 16'd20917, 16'd43274}; // indx = 2495
    #10;
    addra = 32'd79872;
    dina = {96'd0, 16'd47691, 16'd17104, 16'd10346, 16'd54189, 16'd31085, 16'd31302, 16'd51952, 16'd49079, 16'd64421, 16'd25378}; // indx = 2496
    #10;
    addra = 32'd79904;
    dina = {96'd0, 16'd38930, 16'd6521, 16'd12191, 16'd49419, 16'd9272, 16'd65279, 16'd31719, 16'd17668, 16'd21672, 16'd65286}; // indx = 2497
    #10;
    addra = 32'd79936;
    dina = {96'd0, 16'd64132, 16'd61388, 16'd28155, 16'd33110, 16'd12838, 16'd12900, 16'd62728, 16'd17640, 16'd61757, 16'd4206}; // indx = 2498
    #10;
    addra = 32'd79968;
    dina = {96'd0, 16'd62109, 16'd54740, 16'd63228, 16'd64670, 16'd48165, 16'd22337, 16'd65238, 16'd36866, 16'd4910, 16'd63298}; // indx = 2499
    #10;
    addra = 32'd80000;
    dina = {96'd0, 16'd47423, 16'd52208, 16'd41653, 16'd25787, 16'd50635, 16'd17375, 16'd30462, 16'd51398, 16'd38858, 16'd49838}; // indx = 2500
    #10;
    addra = 32'd80032;
    dina = {96'd0, 16'd57799, 16'd15194, 16'd9754, 16'd27287, 16'd50983, 16'd63693, 16'd25849, 16'd5515, 16'd29444, 16'd25497}; // indx = 2501
    #10;
    addra = 32'd80064;
    dina = {96'd0, 16'd17416, 16'd54946, 16'd25598, 16'd37377, 16'd9128, 16'd38840, 16'd41080, 16'd47590, 16'd55915, 16'd58371}; // indx = 2502
    #10;
    addra = 32'd80096;
    dina = {96'd0, 16'd10777, 16'd22309, 16'd49794, 16'd58131, 16'd769, 16'd20766, 16'd63149, 16'd14240, 16'd2210, 16'd44392}; // indx = 2503
    #10;
    addra = 32'd80128;
    dina = {96'd0, 16'd47263, 16'd54695, 16'd12440, 16'd34553, 16'd17136, 16'd29809, 16'd22671, 16'd45051, 16'd30438, 16'd22380}; // indx = 2504
    #10;
    addra = 32'd80160;
    dina = {96'd0, 16'd52064, 16'd61526, 16'd45977, 16'd32397, 16'd49616, 16'd17, 16'd27051, 16'd61452, 16'd65071, 16'd46085}; // indx = 2505
    #10;
    addra = 32'd80192;
    dina = {96'd0, 16'd2182, 16'd51082, 16'd42163, 16'd25381, 16'd10463, 16'd44822, 16'd4444, 16'd55016, 16'd43608, 16'd26402}; // indx = 2506
    #10;
    addra = 32'd80224;
    dina = {96'd0, 16'd35916, 16'd52498, 16'd8046, 16'd28792, 16'd5181, 16'd695, 16'd10170, 16'd42121, 16'd50120, 16'd20859}; // indx = 2507
    #10;
    addra = 32'd80256;
    dina = {96'd0, 16'd17890, 16'd37751, 16'd11848, 16'd54448, 16'd37620, 16'd49868, 16'd31591, 16'd63160, 16'd55453, 16'd22612}; // indx = 2508
    #10;
    addra = 32'd80288;
    dina = {96'd0, 16'd19576, 16'd14366, 16'd22787, 16'd2932, 16'd1589, 16'd61690, 16'd61414, 16'd54636, 16'd64572, 16'd32173}; // indx = 2509
    #10;
    addra = 32'd80320;
    dina = {96'd0, 16'd52568, 16'd36222, 16'd19890, 16'd39878, 16'd7463, 16'd47924, 16'd7098, 16'd6735, 16'd30534, 16'd34271}; // indx = 2510
    #10;
    addra = 32'd80352;
    dina = {96'd0, 16'd42678, 16'd59704, 16'd26256, 16'd7648, 16'd36417, 16'd6066, 16'd25653, 16'd19280, 16'd23558, 16'd55346}; // indx = 2511
    #10;
    addra = 32'd80384;
    dina = {96'd0, 16'd15267, 16'd17855, 16'd50035, 16'd26808, 16'd64184, 16'd33526, 16'd11913, 16'd10922, 16'd30234, 16'd36309}; // indx = 2512
    #10;
    addra = 32'd80416;
    dina = {96'd0, 16'd18821, 16'd52196, 16'd62015, 16'd61957, 16'd21664, 16'd729, 16'd10793, 16'd46036, 16'd16945, 16'd20009}; // indx = 2513
    #10;
    addra = 32'd80448;
    dina = {96'd0, 16'd54287, 16'd7241, 16'd27389, 16'd48860, 16'd51272, 16'd24399, 16'd20941, 16'd44175, 16'd52884, 16'd48616}; // indx = 2514
    #10;
    addra = 32'd80480;
    dina = {96'd0, 16'd46563, 16'd1093, 16'd55687, 16'd58368, 16'd10246, 16'd24709, 16'd7309, 16'd45126, 16'd27543, 16'd52509}; // indx = 2515
    #10;
    addra = 32'd80512;
    dina = {96'd0, 16'd13962, 16'd9379, 16'd24408, 16'd19883, 16'd3453, 16'd30763, 16'd27768, 16'd38880, 16'd29562, 16'd23271}; // indx = 2516
    #10;
    addra = 32'd80544;
    dina = {96'd0, 16'd23089, 16'd43747, 16'd51437, 16'd64133, 16'd17254, 16'd64915, 16'd42746, 16'd42393, 16'd17859, 16'd7230}; // indx = 2517
    #10;
    addra = 32'd80576;
    dina = {96'd0, 16'd13237, 16'd36803, 16'd958, 16'd10981, 16'd55743, 16'd65441, 16'd4819, 16'd40672, 16'd19906, 16'd4645}; // indx = 2518
    #10;
    addra = 32'd80608;
    dina = {96'd0, 16'd56430, 16'd49099, 16'd7807, 16'd9252, 16'd13030, 16'd5539, 16'd62418, 16'd21952, 16'd1558, 16'd18162}; // indx = 2519
    #10;
    addra = 32'd80640;
    dina = {96'd0, 16'd23853, 16'd18970, 16'd26226, 16'd51616, 16'd25882, 16'd35731, 16'd3948, 16'd26135, 16'd31741, 16'd25043}; // indx = 2520
    #10;
    addra = 32'd80672;
    dina = {96'd0, 16'd30357, 16'd49420, 16'd63427, 16'd21484, 16'd28441, 16'd26412, 16'd43970, 16'd13348, 16'd47946, 16'd46571}; // indx = 2521
    #10;
    addra = 32'd80704;
    dina = {96'd0, 16'd26761, 16'd45919, 16'd55491, 16'd62407, 16'd34087, 16'd54130, 16'd21222, 16'd9369, 16'd12576, 16'd57480}; // indx = 2522
    #10;
    addra = 32'd80736;
    dina = {96'd0, 16'd37555, 16'd29402, 16'd11605, 16'd50645, 16'd11382, 16'd33219, 16'd10859, 16'd16465, 16'd13301, 16'd42485}; // indx = 2523
    #10;
    addra = 32'd80768;
    dina = {96'd0, 16'd48762, 16'd17441, 16'd20709, 16'd63696, 16'd11920, 16'd62266, 16'd43423, 16'd45481, 16'd49758, 16'd44893}; // indx = 2524
    #10;
    addra = 32'd80800;
    dina = {96'd0, 16'd43402, 16'd47696, 16'd4242, 16'd50492, 16'd39998, 16'd50509, 16'd13629, 16'd63556, 16'd2846, 16'd16645}; // indx = 2525
    #10;
    addra = 32'd80832;
    dina = {96'd0, 16'd9160, 16'd2558, 16'd51454, 16'd42615, 16'd22629, 16'd29645, 16'd50807, 16'd37430, 16'd57703, 16'd9460}; // indx = 2526
    #10;
    addra = 32'd80864;
    dina = {96'd0, 16'd32793, 16'd28506, 16'd11540, 16'd23562, 16'd32673, 16'd27592, 16'd45922, 16'd28588, 16'd1801, 16'd31344}; // indx = 2527
    #10;
    addra = 32'd80896;
    dina = {96'd0, 16'd44955, 16'd49650, 16'd33637, 16'd44210, 16'd7303, 16'd3459, 16'd55835, 16'd45585, 16'd55276, 16'd7187}; // indx = 2528
    #10;
    addra = 32'd80928;
    dina = {96'd0, 16'd27582, 16'd32293, 16'd25761, 16'd33896, 16'd10877, 16'd3794, 16'd42504, 16'd46259, 16'd26027, 16'd15581}; // indx = 2529
    #10;
    addra = 32'd80960;
    dina = {96'd0, 16'd688, 16'd234, 16'd23277, 16'd52454, 16'd31389, 16'd57196, 16'd34840, 16'd1516, 16'd33646, 16'd35878}; // indx = 2530
    #10;
    addra = 32'd80992;
    dina = {96'd0, 16'd4480, 16'd21209, 16'd35288, 16'd55907, 16'd30726, 16'd14104, 16'd24458, 16'd43717, 16'd60688, 16'd23173}; // indx = 2531
    #10;
    addra = 32'd81024;
    dina = {96'd0, 16'd29053, 16'd13899, 16'd59942, 16'd34665, 16'd49631, 16'd10877, 16'd54361, 16'd28215, 16'd37810, 16'd57287}; // indx = 2532
    #10;
    addra = 32'd81056;
    dina = {96'd0, 16'd31775, 16'd29861, 16'd29065, 16'd11361, 16'd17865, 16'd27987, 16'd25712, 16'd16599, 16'd32398, 16'd15247}; // indx = 2533
    #10;
    addra = 32'd81088;
    dina = {96'd0, 16'd7913, 16'd48237, 16'd49466, 16'd5485, 16'd29345, 16'd26459, 16'd22441, 16'd12555, 16'd16636, 16'd1033}; // indx = 2534
    #10;
    addra = 32'd81120;
    dina = {96'd0, 16'd62324, 16'd11789, 16'd54686, 16'd62962, 16'd8843, 16'd42808, 16'd23571, 16'd4993, 16'd42407, 16'd2787}; // indx = 2535
    #10;
    addra = 32'd81152;
    dina = {96'd0, 16'd36584, 16'd25567, 16'd26894, 16'd9971, 16'd56505, 16'd35477, 16'd61212, 16'd9484, 16'd17305, 16'd60417}; // indx = 2536
    #10;
    addra = 32'd81184;
    dina = {96'd0, 16'd14293, 16'd30027, 16'd7227, 16'd3755, 16'd39993, 16'd65104, 16'd19758, 16'd6518, 16'd47936, 16'd2828}; // indx = 2537
    #10;
    addra = 32'd81216;
    dina = {96'd0, 16'd11154, 16'd25349, 16'd37783, 16'd23634, 16'd26249, 16'd27366, 16'd21102, 16'd23361, 16'd41076, 16'd5980}; // indx = 2538
    #10;
    addra = 32'd81248;
    dina = {96'd0, 16'd31966, 16'd31347, 16'd44422, 16'd40095, 16'd30709, 16'd51440, 16'd16662, 16'd55153, 16'd63080, 16'd29407}; // indx = 2539
    #10;
    addra = 32'd81280;
    dina = {96'd0, 16'd29123, 16'd16088, 16'd53640, 16'd61184, 16'd4807, 16'd28208, 16'd29206, 16'd32064, 16'd2174, 16'd65138}; // indx = 2540
    #10;
    addra = 32'd81312;
    dina = {96'd0, 16'd6436, 16'd9940, 16'd62986, 16'd40203, 16'd19973, 16'd14563, 16'd20790, 16'd54909, 16'd22619, 16'd11999}; // indx = 2541
    #10;
    addra = 32'd81344;
    dina = {96'd0, 16'd34269, 16'd11510, 16'd60063, 16'd58371, 16'd4402, 16'd50592, 16'd10794, 16'd1955, 16'd20120, 16'd45372}; // indx = 2542
    #10;
    addra = 32'd81376;
    dina = {96'd0, 16'd24258, 16'd41656, 16'd35938, 16'd41372, 16'd23037, 16'd31566, 16'd2853, 16'd9906, 16'd34006, 16'd45868}; // indx = 2543
    #10;
    addra = 32'd81408;
    dina = {96'd0, 16'd29471, 16'd50803, 16'd36078, 16'd33996, 16'd11290, 16'd5132, 16'd24508, 16'd10338, 16'd8716, 16'd53303}; // indx = 2544
    #10;
    addra = 32'd81440;
    dina = {96'd0, 16'd22823, 16'd27733, 16'd23914, 16'd12606, 16'd39278, 16'd9587, 16'd48977, 16'd42401, 16'd5003, 16'd19673}; // indx = 2545
    #10;
    addra = 32'd81472;
    dina = {96'd0, 16'd13, 16'd25560, 16'd33049, 16'd65016, 16'd30942, 16'd25856, 16'd14984, 16'd7012, 16'd6072, 16'd53946}; // indx = 2546
    #10;
    addra = 32'd81504;
    dina = {96'd0, 16'd5556, 16'd22095, 16'd52151, 16'd24492, 16'd62073, 16'd10294, 16'd38514, 16'd44531, 16'd38542, 16'd20510}; // indx = 2547
    #10;
    addra = 32'd81536;
    dina = {96'd0, 16'd42289, 16'd35646, 16'd60804, 16'd42155, 16'd14251, 16'd64326, 16'd39303, 16'd55326, 16'd13772, 16'd61522}; // indx = 2548
    #10;
    addra = 32'd81568;
    dina = {96'd0, 16'd60823, 16'd23468, 16'd64422, 16'd58366, 16'd26467, 16'd51507, 16'd925, 16'd60181, 16'd13853, 16'd42816}; // indx = 2549
    #10;
    addra = 32'd81600;
    dina = {96'd0, 16'd35620, 16'd18686, 16'd60898, 16'd13025, 16'd2266, 16'd50789, 16'd22838, 16'd64027, 16'd32869, 16'd53096}; // indx = 2550
    #10;
    addra = 32'd81632;
    dina = {96'd0, 16'd20283, 16'd56805, 16'd31708, 16'd31849, 16'd5230, 16'd58965, 16'd32415, 16'd22174, 16'd64827, 16'd12430}; // indx = 2551
    #10;
    addra = 32'd81664;
    dina = {96'd0, 16'd37824, 16'd13842, 16'd52714, 16'd43712, 16'd29936, 16'd41521, 16'd25138, 16'd8699, 16'd18796, 16'd12443}; // indx = 2552
    #10;
    addra = 32'd81696;
    dina = {96'd0, 16'd48406, 16'd912, 16'd13764, 16'd55892, 16'd56510, 16'd14344, 16'd18963, 16'd60986, 16'd63260, 16'd7518}; // indx = 2553
    #10;
    addra = 32'd81728;
    dina = {96'd0, 16'd47736, 16'd243, 16'd15873, 16'd34358, 16'd41057, 16'd6600, 16'd42676, 16'd53069, 16'd45840, 16'd34827}; // indx = 2554
    #10;
    addra = 32'd81760;
    dina = {96'd0, 16'd59947, 16'd12182, 16'd59354, 16'd422, 16'd37889, 16'd31653, 16'd7402, 16'd49744, 16'd6789, 16'd16234}; // indx = 2555
    #10;
    addra = 32'd81792;
    dina = {96'd0, 16'd61928, 16'd36641, 16'd22524, 16'd10505, 16'd55784, 16'd13333, 16'd46047, 16'd48381, 16'd37456, 16'd53043}; // indx = 2556
    #10;
    addra = 32'd81824;
    dina = {96'd0, 16'd31089, 16'd15131, 16'd50181, 16'd23197, 16'd46382, 16'd13323, 16'd52240, 16'd64652, 16'd19245, 16'd45141}; // indx = 2557
    #10;
    addra = 32'd81856;
    dina = {96'd0, 16'd23114, 16'd63976, 16'd31920, 16'd46342, 16'd58001, 16'd28339, 16'd32666, 16'd63912, 16'd19765, 16'd5163}; // indx = 2558
    #10;
    addra = 32'd81888;
    dina = {96'd0, 16'd14912, 16'd10569, 16'd6390, 16'd16375, 16'd12905, 16'd25239, 16'd49056, 16'd59140, 16'd62080, 16'd60270}; // indx = 2559
    #10;
    addra = 32'd81920;
    dina = {96'd0, 16'd26710, 16'd36354, 16'd18150, 16'd26448, 16'd33758, 16'd5862, 16'd62912, 16'd45942, 16'd14819, 16'd31863}; // indx = 2560
    #10;
    addra = 32'd81952;
    dina = {96'd0, 16'd16502, 16'd51908, 16'd33118, 16'd59738, 16'd40503, 16'd18173, 16'd48935, 16'd40100, 16'd1636, 16'd45302}; // indx = 2561
    #10;
    addra = 32'd81984;
    dina = {96'd0, 16'd58807, 16'd6197, 16'd2970, 16'd26764, 16'd54863, 16'd60326, 16'd54023, 16'd24023, 16'd7119, 16'd57296}; // indx = 2562
    #10;
    addra = 32'd82016;
    dina = {96'd0, 16'd47804, 16'd16421, 16'd451, 16'd34268, 16'd58085, 16'd20371, 16'd5041, 16'd58585, 16'd6711, 16'd22705}; // indx = 2563
    #10;
    addra = 32'd82048;
    dina = {96'd0, 16'd45235, 16'd4624, 16'd43855, 16'd22522, 16'd46380, 16'd9453, 16'd8447, 16'd54022, 16'd55671, 16'd8456}; // indx = 2564
    #10;
    addra = 32'd82080;
    dina = {96'd0, 16'd15199, 16'd5683, 16'd25989, 16'd32503, 16'd57174, 16'd37540, 16'd62144, 16'd18297, 16'd51431, 16'd7678}; // indx = 2565
    #10;
    addra = 32'd82112;
    dina = {96'd0, 16'd52105, 16'd169, 16'd240, 16'd28433, 16'd57127, 16'd20100, 16'd10006, 16'd612, 16'd58186, 16'd34832}; // indx = 2566
    #10;
    addra = 32'd82144;
    dina = {96'd0, 16'd36125, 16'd57382, 16'd8839, 16'd145, 16'd40890, 16'd64261, 16'd35890, 16'd65038, 16'd63169, 16'd62595}; // indx = 2567
    #10;
    addra = 32'd82176;
    dina = {96'd0, 16'd19623, 16'd28685, 16'd48629, 16'd17281, 16'd55941, 16'd21113, 16'd29859, 16'd62775, 16'd50069, 16'd21411}; // indx = 2568
    #10;
    addra = 32'd82208;
    dina = {96'd0, 16'd34134, 16'd7709, 16'd37931, 16'd42107, 16'd3412, 16'd21401, 16'd64777, 16'd18396, 16'd38751, 16'd27217}; // indx = 2569
    #10;
    addra = 32'd82240;
    dina = {96'd0, 16'd35337, 16'd28986, 16'd3882, 16'd49172, 16'd43870, 16'd31640, 16'd7320, 16'd9859, 16'd62369, 16'd50510}; // indx = 2570
    #10;
    addra = 32'd82272;
    dina = {96'd0, 16'd57139, 16'd12655, 16'd14631, 16'd25534, 16'd59636, 16'd38481, 16'd15808, 16'd58350, 16'd24397, 16'd35579}; // indx = 2571
    #10;
    addra = 32'd82304;
    dina = {96'd0, 16'd19558, 16'd57814, 16'd6846, 16'd17265, 16'd55896, 16'd47822, 16'd21848, 16'd38861, 16'd52629, 16'd46753}; // indx = 2572
    #10;
    addra = 32'd82336;
    dina = {96'd0, 16'd46679, 16'd3135, 16'd16187, 16'd9735, 16'd15784, 16'd27695, 16'd4924, 16'd50208, 16'd49480, 16'd46246}; // indx = 2573
    #10;
    addra = 32'd82368;
    dina = {96'd0, 16'd48066, 16'd22493, 16'd20141, 16'd2391, 16'd57400, 16'd65118, 16'd20232, 16'd63722, 16'd39700, 16'd43969}; // indx = 2574
    #10;
    addra = 32'd82400;
    dina = {96'd0, 16'd51722, 16'd14783, 16'd37116, 16'd46739, 16'd28825, 16'd25933, 16'd33444, 16'd63328, 16'd55897, 16'd35403}; // indx = 2575
    #10;
    addra = 32'd82432;
    dina = {96'd0, 16'd55108, 16'd25834, 16'd52886, 16'd10441, 16'd13109, 16'd58610, 16'd15335, 16'd9149, 16'd26089, 16'd16376}; // indx = 2576
    #10;
    addra = 32'd82464;
    dina = {96'd0, 16'd59693, 16'd23746, 16'd8749, 16'd43893, 16'd12121, 16'd54632, 16'd55595, 16'd27499, 16'd21582, 16'd44841}; // indx = 2577
    #10;
    addra = 32'd82496;
    dina = {96'd0, 16'd32923, 16'd49, 16'd57510, 16'd60009, 16'd23057, 16'd46821, 16'd43929, 16'd5433, 16'd37878, 16'd15185}; // indx = 2578
    #10;
    addra = 32'd82528;
    dina = {96'd0, 16'd48110, 16'd13144, 16'd25781, 16'd28979, 16'd19483, 16'd28622, 16'd61424, 16'd24864, 16'd63631, 16'd15023}; // indx = 2579
    #10;
    addra = 32'd82560;
    dina = {96'd0, 16'd33507, 16'd33976, 16'd35251, 16'd19423, 16'd45530, 16'd26564, 16'd22689, 16'd8121, 16'd44692, 16'd21712}; // indx = 2580
    #10;
    addra = 32'd82592;
    dina = {96'd0, 16'd49119, 16'd60858, 16'd52381, 16'd10942, 16'd26218, 16'd25816, 16'd6948, 16'd48412, 16'd30271, 16'd56831}; // indx = 2581
    #10;
    addra = 32'd82624;
    dina = {96'd0, 16'd51060, 16'd62385, 16'd29130, 16'd14851, 16'd31382, 16'd50322, 16'd24382, 16'd61485, 16'd33832, 16'd22628}; // indx = 2582
    #10;
    addra = 32'd82656;
    dina = {96'd0, 16'd1485, 16'd42548, 16'd31159, 16'd4306, 16'd48302, 16'd11599, 16'd15941, 16'd23461, 16'd5921, 16'd42674}; // indx = 2583
    #10;
    addra = 32'd82688;
    dina = {96'd0, 16'd8033, 16'd3287, 16'd18012, 16'd53238, 16'd47900, 16'd36189, 16'd23453, 16'd35970, 16'd45394, 16'd26960}; // indx = 2584
    #10;
    addra = 32'd82720;
    dina = {96'd0, 16'd39224, 16'd19485, 16'd62569, 16'd47805, 16'd13470, 16'd25231, 16'd18063, 16'd2444, 16'd53762, 16'd6973}; // indx = 2585
    #10;
    addra = 32'd82752;
    dina = {96'd0, 16'd42235, 16'd16190, 16'd16982, 16'd10413, 16'd4400, 16'd619, 16'd6605, 16'd46230, 16'd63410, 16'd64727}; // indx = 2586
    #10;
    addra = 32'd82784;
    dina = {96'd0, 16'd62167, 16'd18165, 16'd15787, 16'd39675, 16'd27500, 16'd23440, 16'd4721, 16'd18714, 16'd65431, 16'd4911}; // indx = 2587
    #10;
    addra = 32'd82816;
    dina = {96'd0, 16'd3949, 16'd55984, 16'd50882, 16'd9027, 16'd16476, 16'd47992, 16'd32989, 16'd47323, 16'd53171, 16'd3181}; // indx = 2588
    #10;
    addra = 32'd82848;
    dina = {96'd0, 16'd49978, 16'd20391, 16'd27928, 16'd50982, 16'd6746, 16'd58822, 16'd52204, 16'd38696, 16'd61884, 16'd25923}; // indx = 2589
    #10;
    addra = 32'd82880;
    dina = {96'd0, 16'd55779, 16'd55607, 16'd51182, 16'd26674, 16'd52062, 16'd22900, 16'd48924, 16'd11115, 16'd21785, 16'd11646}; // indx = 2590
    #10;
    addra = 32'd82912;
    dina = {96'd0, 16'd8405, 16'd49341, 16'd26606, 16'd32091, 16'd53944, 16'd404, 16'd8871, 16'd33591, 16'd51495, 16'd33905}; // indx = 2591
    #10;
    addra = 32'd82944;
    dina = {96'd0, 16'd50142, 16'd46167, 16'd35204, 16'd40994, 16'd50525, 16'd53846, 16'd417, 16'd13706, 16'd20908, 16'd17412}; // indx = 2592
    #10;
    addra = 32'd82976;
    dina = {96'd0, 16'd31317, 16'd51108, 16'd23869, 16'd60399, 16'd51708, 16'd41067, 16'd53118, 16'd43468, 16'd23060, 16'd53124}; // indx = 2593
    #10;
    addra = 32'd83008;
    dina = {96'd0, 16'd9964, 16'd2756, 16'd35765, 16'd61621, 16'd62012, 16'd28997, 16'd8196, 16'd48860, 16'd57146, 16'd30947}; // indx = 2594
    #10;
    addra = 32'd83040;
    dina = {96'd0, 16'd26450, 16'd55324, 16'd53539, 16'd45276, 16'd6469, 16'd464, 16'd51127, 16'd29011, 16'd46372, 16'd9018}; // indx = 2595
    #10;
    addra = 32'd83072;
    dina = {96'd0, 16'd56175, 16'd20185, 16'd17524, 16'd12639, 16'd41308, 16'd10255, 16'd63267, 16'd15473, 16'd19110, 16'd2591}; // indx = 2596
    #10;
    addra = 32'd83104;
    dina = {96'd0, 16'd19902, 16'd46109, 16'd12809, 16'd48308, 16'd51522, 16'd41499, 16'd17979, 16'd31874, 16'd10040, 16'd3664}; // indx = 2597
    #10;
    addra = 32'd83136;
    dina = {96'd0, 16'd49075, 16'd8356, 16'd25797, 16'd28623, 16'd64950, 16'd3372, 16'd26006, 16'd38916, 16'd56464, 16'd51905}; // indx = 2598
    #10;
    addra = 32'd83168;
    dina = {96'd0, 16'd50106, 16'd6969, 16'd37388, 16'd40238, 16'd38570, 16'd2050, 16'd55150, 16'd47958, 16'd13808, 16'd26072}; // indx = 2599
    #10;
    addra = 32'd83200;
    dina = {96'd0, 16'd56702, 16'd40057, 16'd50963, 16'd28528, 16'd27605, 16'd53184, 16'd36858, 16'd31255, 16'd50017, 16'd15933}; // indx = 2600
    #10;
    addra = 32'd83232;
    dina = {96'd0, 16'd12062, 16'd44345, 16'd29574, 16'd22108, 16'd3851, 16'd28916, 16'd7720, 16'd43609, 16'd64557, 16'd27853}; // indx = 2601
    #10;
    addra = 32'd83264;
    dina = {96'd0, 16'd40266, 16'd43962, 16'd58781, 16'd5934, 16'd2895, 16'd29369, 16'd22413, 16'd20263, 16'd32376, 16'd40019}; // indx = 2602
    #10;
    addra = 32'd83296;
    dina = {96'd0, 16'd64149, 16'd21362, 16'd38977, 16'd58067, 16'd9044, 16'd28113, 16'd57863, 16'd61795, 16'd12376, 16'd1008}; // indx = 2603
    #10;
    addra = 32'd83328;
    dina = {96'd0, 16'd5184, 16'd3768, 16'd5860, 16'd16686, 16'd3229, 16'd55092, 16'd62974, 16'd23833, 16'd52972, 16'd61219}; // indx = 2604
    #10;
    addra = 32'd83360;
    dina = {96'd0, 16'd17895, 16'd51237, 16'd43221, 16'd33565, 16'd38154, 16'd13103, 16'd39907, 16'd12330, 16'd58836, 16'd48002}; // indx = 2605
    #10;
    addra = 32'd83392;
    dina = {96'd0, 16'd21302, 16'd3468, 16'd62905, 16'd20800, 16'd9408, 16'd34907, 16'd340, 16'd31543, 16'd18345, 16'd17482}; // indx = 2606
    #10;
    addra = 32'd83424;
    dina = {96'd0, 16'd28636, 16'd39444, 16'd46577, 16'd6198, 16'd16916, 16'd15007, 16'd31714, 16'd18305, 16'd40993, 16'd15688}; // indx = 2607
    #10;
    addra = 32'd83456;
    dina = {96'd0, 16'd37788, 16'd1255, 16'd59833, 16'd13238, 16'd27187, 16'd49566, 16'd38061, 16'd55130, 16'd12161, 16'd40259}; // indx = 2608
    #10;
    addra = 32'd83488;
    dina = {96'd0, 16'd49281, 16'd29337, 16'd21862, 16'd30156, 16'd34377, 16'd23098, 16'd2752, 16'd30347, 16'd30843, 16'd36569}; // indx = 2609
    #10;
    addra = 32'd83520;
    dina = {96'd0, 16'd26017, 16'd22543, 16'd46372, 16'd1779, 16'd17570, 16'd63810, 16'd41489, 16'd56128, 16'd11429, 16'd59584}; // indx = 2610
    #10;
    addra = 32'd83552;
    dina = {96'd0, 16'd13982, 16'd47834, 16'd53211, 16'd29511, 16'd34920, 16'd16714, 16'd65525, 16'd61676, 16'd46449, 16'd10997}; // indx = 2611
    #10;
    addra = 32'd83584;
    dina = {96'd0, 16'd25306, 16'd15944, 16'd10640, 16'd10896, 16'd3429, 16'd36025, 16'd26947, 16'd5022, 16'd11916, 16'd52708}; // indx = 2612
    #10;
    addra = 32'd83616;
    dina = {96'd0, 16'd63259, 16'd20557, 16'd48564, 16'd44749, 16'd5083, 16'd53546, 16'd21779, 16'd1905, 16'd9597, 16'd63609}; // indx = 2613
    #10;
    addra = 32'd83648;
    dina = {96'd0, 16'd32761, 16'd25367, 16'd10074, 16'd41088, 16'd22794, 16'd2794, 16'd46194, 16'd45977, 16'd46379, 16'd11965}; // indx = 2614
    #10;
    addra = 32'd83680;
    dina = {96'd0, 16'd54716, 16'd43236, 16'd25051, 16'd11142, 16'd21893, 16'd48190, 16'd61211, 16'd62420, 16'd18970, 16'd6376}; // indx = 2615
    #10;
    addra = 32'd83712;
    dina = {96'd0, 16'd57257, 16'd36560, 16'd37791, 16'd32855, 16'd24016, 16'd38203, 16'd4944, 16'd45110, 16'd7598, 16'd17689}; // indx = 2616
    #10;
    addra = 32'd83744;
    dina = {96'd0, 16'd63745, 16'd63170, 16'd54382, 16'd19639, 16'd42367, 16'd35034, 16'd15558, 16'd15314, 16'd31397, 16'd29437}; // indx = 2617
    #10;
    addra = 32'd83776;
    dina = {96'd0, 16'd15910, 16'd48411, 16'd43426, 16'd60285, 16'd25698, 16'd6593, 16'd40549, 16'd9428, 16'd4708, 16'd2285}; // indx = 2618
    #10;
    addra = 32'd83808;
    dina = {96'd0, 16'd27848, 16'd43982, 16'd31615, 16'd39943, 16'd61897, 16'd2500, 16'd62954, 16'd11711, 16'd43551, 16'd29818}; // indx = 2619
    #10;
    addra = 32'd83840;
    dina = {96'd0, 16'd42354, 16'd64512, 16'd41359, 16'd14235, 16'd60660, 16'd30526, 16'd59872, 16'd39466, 16'd25781, 16'd38004}; // indx = 2620
    #10;
    addra = 32'd83872;
    dina = {96'd0, 16'd39714, 16'd41323, 16'd34436, 16'd33115, 16'd11827, 16'd22367, 16'd42388, 16'd1164, 16'd18798, 16'd59464}; // indx = 2621
    #10;
    addra = 32'd83904;
    dina = {96'd0, 16'd9424, 16'd46366, 16'd48247, 16'd31235, 16'd1037, 16'd59774, 16'd41579, 16'd51803, 16'd36979, 16'd10571}; // indx = 2622
    #10;
    addra = 32'd83936;
    dina = {96'd0, 16'd2565, 16'd6183, 16'd8276, 16'd1244, 16'd54576, 16'd3386, 16'd63839, 16'd4237, 16'd61708, 16'd52423}; // indx = 2623
    #10;
    addra = 32'd83968;
    dina = {96'd0, 16'd6109, 16'd10847, 16'd26983, 16'd4785, 16'd56377, 16'd51590, 16'd1693, 16'd21217, 16'd26574, 16'd10634}; // indx = 2624
    #10;
    addra = 32'd84000;
    dina = {96'd0, 16'd35046, 16'd6829, 16'd17993, 16'd23433, 16'd43263, 16'd5232, 16'd52616, 16'd24441, 16'd25413, 16'd25965}; // indx = 2625
    #10;
    addra = 32'd84032;
    dina = {96'd0, 16'd57230, 16'd57335, 16'd45878, 16'd59544, 16'd16666, 16'd38644, 16'd57907, 16'd33501, 16'd34505, 16'd18133}; // indx = 2626
    #10;
    addra = 32'd84064;
    dina = {96'd0, 16'd58642, 16'd55195, 16'd61357, 16'd41965, 16'd40802, 16'd46664, 16'd17581, 16'd58604, 16'd21245, 16'd21898}; // indx = 2627
    #10;
    addra = 32'd84096;
    dina = {96'd0, 16'd29872, 16'd33949, 16'd4410, 16'd15035, 16'd89, 16'd57272, 16'd17158, 16'd22036, 16'd6752, 16'd22621}; // indx = 2628
    #10;
    addra = 32'd84128;
    dina = {96'd0, 16'd43299, 16'd43232, 16'd17433, 16'd18728, 16'd41220, 16'd56591, 16'd7247, 16'd39128, 16'd62102, 16'd36542}; // indx = 2629
    #10;
    addra = 32'd84160;
    dina = {96'd0, 16'd44862, 16'd64471, 16'd42849, 16'd58204, 16'd38967, 16'd16947, 16'd61655, 16'd30718, 16'd61717, 16'd35725}; // indx = 2630
    #10;
    addra = 32'd84192;
    dina = {96'd0, 16'd23249, 16'd4411, 16'd42787, 16'd18956, 16'd4042, 16'd51392, 16'd11381, 16'd9506, 16'd9246, 16'd18796}; // indx = 2631
    #10;
    addra = 32'd84224;
    dina = {96'd0, 16'd37587, 16'd17201, 16'd62129, 16'd9129, 16'd21873, 16'd62834, 16'd17349, 16'd25807, 16'd13693, 16'd41349}; // indx = 2632
    #10;
    addra = 32'd84256;
    dina = {96'd0, 16'd60790, 16'd49070, 16'd37084, 16'd51427, 16'd56145, 16'd49504, 16'd21412, 16'd33719, 16'd62761, 16'd43171}; // indx = 2633
    #10;
    addra = 32'd84288;
    dina = {96'd0, 16'd47212, 16'd38501, 16'd20389, 16'd2634, 16'd56180, 16'd36173, 16'd56312, 16'd57985, 16'd9616, 16'd36821}; // indx = 2634
    #10;
    addra = 32'd84320;
    dina = {96'd0, 16'd36394, 16'd28239, 16'd1050, 16'd38135, 16'd51346, 16'd43889, 16'd37439, 16'd6581, 16'd35187, 16'd25231}; // indx = 2635
    #10;
    addra = 32'd84352;
    dina = {96'd0, 16'd35301, 16'd889, 16'd224, 16'd32404, 16'd35660, 16'd4068, 16'd32450, 16'd20826, 16'd57421, 16'd44499}; // indx = 2636
    #10;
    addra = 32'd84384;
    dina = {96'd0, 16'd37950, 16'd19974, 16'd27761, 16'd60393, 16'd12648, 16'd1876, 16'd10175, 16'd17477, 16'd38768, 16'd13229}; // indx = 2637
    #10;
    addra = 32'd84416;
    dina = {96'd0, 16'd32171, 16'd24182, 16'd30176, 16'd14075, 16'd48272, 16'd59944, 16'd5495, 16'd41651, 16'd47209, 16'd3971}; // indx = 2638
    #10;
    addra = 32'd84448;
    dina = {96'd0, 16'd12976, 16'd10909, 16'd50031, 16'd40538, 16'd3420, 16'd33823, 16'd18092, 16'd35832, 16'd24613, 16'd61299}; // indx = 2639
    #10;
    addra = 32'd84480;
    dina = {96'd0, 16'd46472, 16'd7070, 16'd42232, 16'd44701, 16'd35486, 16'd29825, 16'd64522, 16'd32991, 16'd29207, 16'd55637}; // indx = 2640
    #10;
    addra = 32'd84512;
    dina = {96'd0, 16'd24606, 16'd32496, 16'd34572, 16'd9811, 16'd24302, 16'd2443, 16'd34332, 16'd21236, 16'd6998, 16'd14568}; // indx = 2641
    #10;
    addra = 32'd84544;
    dina = {96'd0, 16'd63500, 16'd13962, 16'd29058, 16'd8363, 16'd61463, 16'd51853, 16'd17423, 16'd20888, 16'd64143, 16'd46507}; // indx = 2642
    #10;
    addra = 32'd84576;
    dina = {96'd0, 16'd33979, 16'd49907, 16'd60250, 16'd42297, 16'd4137, 16'd43800, 16'd42996, 16'd2061, 16'd29722, 16'd18144}; // indx = 2643
    #10;
    addra = 32'd84608;
    dina = {96'd0, 16'd39923, 16'd56944, 16'd14887, 16'd13129, 16'd1945, 16'd15655, 16'd58074, 16'd53102, 16'd43437, 16'd30799}; // indx = 2644
    #10;
    addra = 32'd84640;
    dina = {96'd0, 16'd57760, 16'd10011, 16'd52676, 16'd56633, 16'd17132, 16'd6193, 16'd10146, 16'd7834, 16'd40097, 16'd6059}; // indx = 2645
    #10;
    addra = 32'd84672;
    dina = {96'd0, 16'd53798, 16'd64269, 16'd44280, 16'd37788, 16'd30932, 16'd20523, 16'd8851, 16'd30098, 16'd3384, 16'd11897}; // indx = 2646
    #10;
    addra = 32'd84704;
    dina = {96'd0, 16'd9907, 16'd7191, 16'd58072, 16'd62718, 16'd9403, 16'd59533, 16'd4164, 16'd41693, 16'd8899, 16'd32094}; // indx = 2647
    #10;
    addra = 32'd84736;
    dina = {96'd0, 16'd5335, 16'd42549, 16'd58696, 16'd16698, 16'd20891, 16'd15718, 16'd35482, 16'd58312, 16'd58246, 16'd43888}; // indx = 2648
    #10;
    addra = 32'd84768;
    dina = {96'd0, 16'd9099, 16'd26205, 16'd33844, 16'd24530, 16'd19536, 16'd24133, 16'd34674, 16'd40410, 16'd3915, 16'd27407}; // indx = 2649
    #10;
    addra = 32'd84800;
    dina = {96'd0, 16'd60787, 16'd23738, 16'd62167, 16'd31711, 16'd20324, 16'd60177, 16'd62363, 16'd36295, 16'd54637, 16'd60834}; // indx = 2650
    #10;
    addra = 32'd84832;
    dina = {96'd0, 16'd50418, 16'd40, 16'd49254, 16'd51874, 16'd12297, 16'd19556, 16'd38813, 16'd2172, 16'd33378, 16'd11663}; // indx = 2651
    #10;
    addra = 32'd84864;
    dina = {96'd0, 16'd34994, 16'd59000, 16'd57210, 16'd54349, 16'd30479, 16'd33513, 16'd52727, 16'd52421, 16'd47046, 16'd43731}; // indx = 2652
    #10;
    addra = 32'd84896;
    dina = {96'd0, 16'd62824, 16'd7299, 16'd13422, 16'd7225, 16'd37145, 16'd22213, 16'd1874, 16'd62516, 16'd3026, 16'd40438}; // indx = 2653
    #10;
    addra = 32'd84928;
    dina = {96'd0, 16'd10297, 16'd7094, 16'd55493, 16'd5410, 16'd21723, 16'd63100, 16'd5667, 16'd35278, 16'd2607, 16'd58111}; // indx = 2654
    #10;
    addra = 32'd84960;
    dina = {96'd0, 16'd47821, 16'd34874, 16'd24403, 16'd23844, 16'd65535, 16'd3836, 16'd52083, 16'd20467, 16'd13447, 16'd20877}; // indx = 2655
    #10;
    addra = 32'd84992;
    dina = {96'd0, 16'd23182, 16'd51398, 16'd47520, 16'd51423, 16'd13732, 16'd4192, 16'd48414, 16'd24649, 16'd31280, 16'd12175}; // indx = 2656
    #10;
    addra = 32'd85024;
    dina = {96'd0, 16'd26454, 16'd22165, 16'd23736, 16'd6390, 16'd52792, 16'd38646, 16'd34070, 16'd13758, 16'd24644, 16'd65185}; // indx = 2657
    #10;
    addra = 32'd85056;
    dina = {96'd0, 16'd21198, 16'd63494, 16'd3959, 16'd50840, 16'd5983, 16'd26198, 16'd64666, 16'd48468, 16'd30433, 16'd64824}; // indx = 2658
    #10;
    addra = 32'd85088;
    dina = {96'd0, 16'd83, 16'd50883, 16'd39308, 16'd47767, 16'd57830, 16'd51788, 16'd36941, 16'd35704, 16'd54916, 16'd58645}; // indx = 2659
    #10;
    addra = 32'd85120;
    dina = {96'd0, 16'd44256, 16'd54302, 16'd37819, 16'd14497, 16'd61096, 16'd55268, 16'd11785, 16'd6368, 16'd64220, 16'd50688}; // indx = 2660
    #10;
    addra = 32'd85152;
    dina = {96'd0, 16'd19109, 16'd49025, 16'd50394, 16'd44411, 16'd6398, 16'd46981, 16'd4496, 16'd26685, 16'd33586, 16'd47962}; // indx = 2661
    #10;
    addra = 32'd85184;
    dina = {96'd0, 16'd7184, 16'd23993, 16'd7451, 16'd26054, 16'd5479, 16'd60441, 16'd49163, 16'd21772, 16'd15599, 16'd27386}; // indx = 2662
    #10;
    addra = 32'd85216;
    dina = {96'd0, 16'd62160, 16'd16247, 16'd52515, 16'd42506, 16'd39408, 16'd24882, 16'd20695, 16'd586, 16'd13203, 16'd19895}; // indx = 2663
    #10;
    addra = 32'd85248;
    dina = {96'd0, 16'd20037, 16'd52047, 16'd36781, 16'd47025, 16'd25271, 16'd30995, 16'd55045, 16'd31253, 16'd7103, 16'd6304}; // indx = 2664
    #10;
    addra = 32'd85280;
    dina = {96'd0, 16'd29987, 16'd10005, 16'd62430, 16'd39650, 16'd49875, 16'd57652, 16'd29866, 16'd23184, 16'd37499, 16'd26353}; // indx = 2665
    #10;
    addra = 32'd85312;
    dina = {96'd0, 16'd18306, 16'd23486, 16'd51644, 16'd18932, 16'd21832, 16'd1016, 16'd51190, 16'd6159, 16'd31343, 16'd9299}; // indx = 2666
    #10;
    addra = 32'd85344;
    dina = {96'd0, 16'd28692, 16'd2190, 16'd52305, 16'd36290, 16'd44117, 16'd11041, 16'd11999, 16'd6962, 16'd32905, 16'd41819}; // indx = 2667
    #10;
    addra = 32'd85376;
    dina = {96'd0, 16'd23191, 16'd54079, 16'd13250, 16'd10100, 16'd27141, 16'd49882, 16'd56749, 16'd44069, 16'd51945, 16'd59456}; // indx = 2668
    #10;
    addra = 32'd85408;
    dina = {96'd0, 16'd14841, 16'd54203, 16'd60728, 16'd20738, 16'd21295, 16'd12980, 16'd56164, 16'd45498, 16'd20693, 16'd25662}; // indx = 2669
    #10;
    addra = 32'd85440;
    dina = {96'd0, 16'd39391, 16'd62257, 16'd65250, 16'd6790, 16'd62551, 16'd7573, 16'd62646, 16'd10519, 16'd57320, 16'd33379}; // indx = 2670
    #10;
    addra = 32'd85472;
    dina = {96'd0, 16'd50286, 16'd28156, 16'd38198, 16'd32364, 16'd55132, 16'd63102, 16'd62787, 16'd15292, 16'd62250, 16'd10137}; // indx = 2671
    #10;
    addra = 32'd85504;
    dina = {96'd0, 16'd6843, 16'd50373, 16'd9074, 16'd39819, 16'd32217, 16'd64250, 16'd21881, 16'd21983, 16'd43983, 16'd60926}; // indx = 2672
    #10;
    addra = 32'd85536;
    dina = {96'd0, 16'd41231, 16'd2433, 16'd54889, 16'd35942, 16'd55408, 16'd42753, 16'd62813, 16'd36861, 16'd49396, 16'd15152}; // indx = 2673
    #10;
    addra = 32'd85568;
    dina = {96'd0, 16'd51717, 16'd13766, 16'd35585, 16'd15156, 16'd65239, 16'd6226, 16'd8237, 16'd28649, 16'd56967, 16'd25203}; // indx = 2674
    #10;
    addra = 32'd85600;
    dina = {96'd0, 16'd49847, 16'd64501, 16'd63155, 16'd38967, 16'd23673, 16'd37507, 16'd63915, 16'd33313, 16'd64731, 16'd34654}; // indx = 2675
    #10;
    addra = 32'd85632;
    dina = {96'd0, 16'd21354, 16'd62840, 16'd33428, 16'd29737, 16'd22584, 16'd5085, 16'd9358, 16'd51823, 16'd34518, 16'd26224}; // indx = 2676
    #10;
    addra = 32'd85664;
    dina = {96'd0, 16'd22384, 16'd65229, 16'd60542, 16'd62516, 16'd18857, 16'd60422, 16'd49887, 16'd65377, 16'd52507, 16'd40576}; // indx = 2677
    #10;
    addra = 32'd85696;
    dina = {96'd0, 16'd12734, 16'd16054, 16'd47822, 16'd34913, 16'd37, 16'd27513, 16'd46424, 16'd54370, 16'd35741, 16'd15595}; // indx = 2678
    #10;
    addra = 32'd85728;
    dina = {96'd0, 16'd15592, 16'd39991, 16'd52862, 16'd59179, 16'd41939, 16'd11049, 16'd12971, 16'd47822, 16'd39700, 16'd3658}; // indx = 2679
    #10;
    addra = 32'd85760;
    dina = {96'd0, 16'd18962, 16'd52108, 16'd53896, 16'd7304, 16'd59602, 16'd31498, 16'd16618, 16'd43130, 16'd47870, 16'd59819}; // indx = 2680
    #10;
    addra = 32'd85792;
    dina = {96'd0, 16'd19018, 16'd42038, 16'd16325, 16'd47818, 16'd56591, 16'd19875, 16'd57727, 16'd63115, 16'd13819, 16'd28079}; // indx = 2681
    #10;
    addra = 32'd85824;
    dina = {96'd0, 16'd35095, 16'd25551, 16'd13626, 16'd29029, 16'd52959, 16'd11440, 16'd46873, 16'd52766, 16'd9495, 16'd2393}; // indx = 2682
    #10;
    addra = 32'd85856;
    dina = {96'd0, 16'd61850, 16'd58528, 16'd42572, 16'd63082, 16'd1873, 16'd26936, 16'd28734, 16'd16286, 16'd54405, 16'd25365}; // indx = 2683
    #10;
    addra = 32'd85888;
    dina = {96'd0, 16'd34440, 16'd34157, 16'd65499, 16'd20662, 16'd38770, 16'd2238, 16'd20322, 16'd44679, 16'd49605, 16'd44461}; // indx = 2684
    #10;
    addra = 32'd85920;
    dina = {96'd0, 16'd2259, 16'd40997, 16'd14813, 16'd21950, 16'd17661, 16'd44929, 16'd39074, 16'd45002, 16'd5280, 16'd47696}; // indx = 2685
    #10;
    addra = 32'd85952;
    dina = {96'd0, 16'd58790, 16'd62195, 16'd41022, 16'd630, 16'd51614, 16'd52478, 16'd61842, 16'd41919, 16'd62385, 16'd18211}; // indx = 2686
    #10;
    addra = 32'd85984;
    dina = {96'd0, 16'd40487, 16'd29741, 16'd13491, 16'd58470, 16'd36758, 16'd33476, 16'd58337, 16'd16848, 16'd30957, 16'd26124}; // indx = 2687
    #10;
    addra = 32'd86016;
    dina = {96'd0, 16'd47098, 16'd40981, 16'd23086, 16'd28349, 16'd44819, 16'd20319, 16'd7316, 16'd17260, 16'd26168, 16'd47543}; // indx = 2688
    #10;
    addra = 32'd86048;
    dina = {96'd0, 16'd51956, 16'd62224, 16'd43321, 16'd39084, 16'd47982, 16'd48605, 16'd63822, 16'd55388, 16'd15963, 16'd27000}; // indx = 2689
    #10;
    addra = 32'd86080;
    dina = {96'd0, 16'd2021, 16'd15319, 16'd26980, 16'd31576, 16'd56350, 16'd16022, 16'd15253, 16'd39122, 16'd7257, 16'd9391}; // indx = 2690
    #10;
    addra = 32'd86112;
    dina = {96'd0, 16'd59287, 16'd42482, 16'd50560, 16'd12272, 16'd50788, 16'd3643, 16'd51985, 16'd30550, 16'd58508, 16'd50419}; // indx = 2691
    #10;
    addra = 32'd86144;
    dina = {96'd0, 16'd17856, 16'd43665, 16'd58719, 16'd42017, 16'd27877, 16'd40039, 16'd36628, 16'd18766, 16'd58883, 16'd35712}; // indx = 2692
    #10;
    addra = 32'd86176;
    dina = {96'd0, 16'd46598, 16'd15530, 16'd32839, 16'd41889, 16'd62450, 16'd11595, 16'd54967, 16'd37213, 16'd702, 16'd53792}; // indx = 2693
    #10;
    addra = 32'd86208;
    dina = {96'd0, 16'd29380, 16'd979, 16'd42052, 16'd9692, 16'd17178, 16'd16011, 16'd18712, 16'd14718, 16'd22559, 16'd50782}; // indx = 2694
    #10;
    addra = 32'd86240;
    dina = {96'd0, 16'd11600, 16'd26102, 16'd9942, 16'd44355, 16'd33851, 16'd49870, 16'd43888, 16'd65078, 16'd42817, 16'd64838}; // indx = 2695
    #10;
    addra = 32'd86272;
    dina = {96'd0, 16'd58568, 16'd5372, 16'd30985, 16'd56666, 16'd43078, 16'd13767, 16'd24374, 16'd17630, 16'd6841, 16'd43721}; // indx = 2696
    #10;
    addra = 32'd86304;
    dina = {96'd0, 16'd62130, 16'd9587, 16'd55687, 16'd28200, 16'd11325, 16'd5968, 16'd7572, 16'd34783, 16'd55120, 16'd48326}; // indx = 2697
    #10;
    addra = 32'd86336;
    dina = {96'd0, 16'd21341, 16'd13036, 16'd56886, 16'd37714, 16'd29318, 16'd31811, 16'd26222, 16'd44607, 16'd20016, 16'd16846}; // indx = 2698
    #10;
    addra = 32'd86368;
    dina = {96'd0, 16'd44207, 16'd27509, 16'd43033, 16'd6847, 16'd45027, 16'd33847, 16'd52371, 16'd44635, 16'd61422, 16'd2772}; // indx = 2699
    #10;
    addra = 32'd86400;
    dina = {96'd0, 16'd30190, 16'd56509, 16'd50586, 16'd18856, 16'd28203, 16'd52970, 16'd50589, 16'd60954, 16'd18179, 16'd60748}; // indx = 2700
    #10;
    addra = 32'd86432;
    dina = {96'd0, 16'd16549, 16'd46094, 16'd21479, 16'd42944, 16'd973, 16'd7514, 16'd57759, 16'd58528, 16'd52471, 16'd33221}; // indx = 2701
    #10;
    addra = 32'd86464;
    dina = {96'd0, 16'd3089, 16'd50226, 16'd57277, 16'd49428, 16'd62078, 16'd42390, 16'd10424, 16'd34966, 16'd46294, 16'd45867}; // indx = 2702
    #10;
    addra = 32'd86496;
    dina = {96'd0, 16'd15030, 16'd30682, 16'd15681, 16'd11922, 16'd25074, 16'd16416, 16'd6763, 16'd34738, 16'd57341, 16'd32662}; // indx = 2703
    #10;
    addra = 32'd86528;
    dina = {96'd0, 16'd57725, 16'd10738, 16'd20778, 16'd64746, 16'd54639, 16'd60021, 16'd86, 16'd18512, 16'd49845, 16'd21490}; // indx = 2704
    #10;
    addra = 32'd86560;
    dina = {96'd0, 16'd4463, 16'd11735, 16'd5399, 16'd19504, 16'd17131, 16'd37156, 16'd63593, 16'd4454, 16'd36937, 16'd62500}; // indx = 2705
    #10;
    addra = 32'd86592;
    dina = {96'd0, 16'd7104, 16'd435, 16'd10864, 16'd18957, 16'd18552, 16'd26493, 16'd36161, 16'd65503, 16'd36632, 16'd24322}; // indx = 2706
    #10;
    addra = 32'd86624;
    dina = {96'd0, 16'd35346, 16'd1350, 16'd46530, 16'd50228, 16'd11166, 16'd47851, 16'd38008, 16'd7389, 16'd54312, 16'd31389}; // indx = 2707
    #10;
    addra = 32'd86656;
    dina = {96'd0, 16'd49800, 16'd14103, 16'd6767, 16'd56965, 16'd29200, 16'd39075, 16'd35769, 16'd14552, 16'd17843, 16'd22265}; // indx = 2708
    #10;
    addra = 32'd86688;
    dina = {96'd0, 16'd56301, 16'd30722, 16'd418, 16'd49087, 16'd41967, 16'd15267, 16'd15845, 16'd40291, 16'd55377, 16'd15035}; // indx = 2709
    #10;
    addra = 32'd86720;
    dina = {96'd0, 16'd22116, 16'd26285, 16'd49829, 16'd43093, 16'd20373, 16'd6567, 16'd32333, 16'd47465, 16'd26202, 16'd31439}; // indx = 2710
    #10;
    addra = 32'd86752;
    dina = {96'd0, 16'd8555, 16'd32673, 16'd18706, 16'd51738, 16'd51581, 16'd59556, 16'd29903, 16'd16290, 16'd46325, 16'd22802}; // indx = 2711
    #10;
    addra = 32'd86784;
    dina = {96'd0, 16'd15128, 16'd1168, 16'd34971, 16'd8542, 16'd1853, 16'd33829, 16'd19943, 16'd22951, 16'd64081, 16'd1779}; // indx = 2712
    #10;
    addra = 32'd86816;
    dina = {96'd0, 16'd8102, 16'd2799, 16'd17802, 16'd43967, 16'd42954, 16'd11835, 16'd46626, 16'd8269, 16'd56438, 16'd8645}; // indx = 2713
    #10;
    addra = 32'd86848;
    dina = {96'd0, 16'd40653, 16'd44100, 16'd10579, 16'd63872, 16'd41854, 16'd3795, 16'd64807, 16'd36213, 16'd16380, 16'd27419}; // indx = 2714
    #10;
    addra = 32'd86880;
    dina = {96'd0, 16'd19845, 16'd18355, 16'd41985, 16'd43830, 16'd22692, 16'd51918, 16'd22981, 16'd48773, 16'd31531, 16'd37370}; // indx = 2715
    #10;
    addra = 32'd86912;
    dina = {96'd0, 16'd41997, 16'd49268, 16'd13939, 16'd54535, 16'd49561, 16'd64307, 16'd38891, 16'd60013, 16'd14589, 16'd64898}; // indx = 2716
    #10;
    addra = 32'd86944;
    dina = {96'd0, 16'd47759, 16'd26343, 16'd45293, 16'd365, 16'd4033, 16'd59258, 16'd980, 16'd30601, 16'd23599, 16'd57648}; // indx = 2717
    #10;
    addra = 32'd86976;
    dina = {96'd0, 16'd2252, 16'd47223, 16'd34737, 16'd19499, 16'd31485, 16'd25964, 16'd47285, 16'd38813, 16'd37456, 16'd12241}; // indx = 2718
    #10;
    addra = 32'd87008;
    dina = {96'd0, 16'd61671, 16'd32944, 16'd58380, 16'd60236, 16'd13734, 16'd25566, 16'd41577, 16'd42087, 16'd38232, 16'd44136}; // indx = 2719
    #10;
    addra = 32'd87040;
    dina = {96'd0, 16'd11263, 16'd17155, 16'd11871, 16'd65377, 16'd65157, 16'd17004, 16'd11903, 16'd7441, 16'd56337, 16'd29377}; // indx = 2720
    #10;
    addra = 32'd87072;
    dina = {96'd0, 16'd5798, 16'd30090, 16'd29333, 16'd21822, 16'd22835, 16'd39778, 16'd47573, 16'd7029, 16'd46614, 16'd5469}; // indx = 2721
    #10;
    addra = 32'd87104;
    dina = {96'd0, 16'd30003, 16'd61020, 16'd39455, 16'd40654, 16'd13774, 16'd57574, 16'd39932, 16'd23401, 16'd9798, 16'd63423}; // indx = 2722
    #10;
    addra = 32'd87136;
    dina = {96'd0, 16'd19469, 16'd44496, 16'd50117, 16'd54879, 16'd22618, 16'd64997, 16'd6176, 16'd8565, 16'd21798, 16'd37797}; // indx = 2723
    #10;
    addra = 32'd87168;
    dina = {96'd0, 16'd28736, 16'd31522, 16'd61087, 16'd60478, 16'd36970, 16'd24232, 16'd5503, 16'd8733, 16'd31039, 16'd36888}; // indx = 2724
    #10;
    addra = 32'd87200;
    dina = {96'd0, 16'd16730, 16'd19615, 16'd45270, 16'd4121, 16'd39239, 16'd19479, 16'd21220, 16'd30625, 16'd38073, 16'd39851}; // indx = 2725
    #10;
    addra = 32'd87232;
    dina = {96'd0, 16'd33799, 16'd37844, 16'd12636, 16'd51645, 16'd37064, 16'd61529, 16'd49113, 16'd31646, 16'd23065, 16'd21776}; // indx = 2726
    #10;
    addra = 32'd87264;
    dina = {96'd0, 16'd19021, 16'd34497, 16'd44073, 16'd47384, 16'd21300, 16'd21105, 16'd53398, 16'd27983, 16'd2495, 16'd31186}; // indx = 2727
    #10;
    addra = 32'd87296;
    dina = {96'd0, 16'd4832, 16'd63767, 16'd61272, 16'd1153, 16'd63262, 16'd41329, 16'd58633, 16'd32058, 16'd56612, 16'd19277}; // indx = 2728
    #10;
    addra = 32'd87328;
    dina = {96'd0, 16'd36994, 16'd10167, 16'd7542, 16'd1485, 16'd10417, 16'd556, 16'd6357, 16'd58221, 16'd34283, 16'd9606}; // indx = 2729
    #10;
    addra = 32'd87360;
    dina = {96'd0, 16'd22725, 16'd11459, 16'd10030, 16'd35435, 16'd61047, 16'd20729, 16'd56209, 16'd39798, 16'd33720, 16'd5737}; // indx = 2730
    #10;
    addra = 32'd87392;
    dina = {96'd0, 16'd60045, 16'd43499, 16'd11297, 16'd14592, 16'd7244, 16'd48149, 16'd45957, 16'd19614, 16'd21035, 16'd36088}; // indx = 2731
    #10;
    addra = 32'd87424;
    dina = {96'd0, 16'd7908, 16'd5691, 16'd26905, 16'd31061, 16'd31550, 16'd40993, 16'd55483, 16'd43116, 16'd6173, 16'd36532}; // indx = 2732
    #10;
    addra = 32'd87456;
    dina = {96'd0, 16'd44766, 16'd58633, 16'd26481, 16'd34048, 16'd39844, 16'd51328, 16'd47815, 16'd31840, 16'd46714, 16'd32779}; // indx = 2733
    #10;
    addra = 32'd87488;
    dina = {96'd0, 16'd39763, 16'd14820, 16'd34678, 16'd50253, 16'd19368, 16'd30430, 16'd11918, 16'd64013, 16'd57879, 16'd19041}; // indx = 2734
    #10;
    addra = 32'd87520;
    dina = {96'd0, 16'd48009, 16'd5265, 16'd49495, 16'd35870, 16'd59414, 16'd12091, 16'd56581, 16'd28986, 16'd35026, 16'd63603}; // indx = 2735
    #10;
    addra = 32'd87552;
    dina = {96'd0, 16'd23227, 16'd49435, 16'd9848, 16'd7430, 16'd43250, 16'd22629, 16'd32519, 16'd19085, 16'd5527, 16'd49577}; // indx = 2736
    #10;
    addra = 32'd87584;
    dina = {96'd0, 16'd62373, 16'd11875, 16'd62255, 16'd30661, 16'd42102, 16'd42558, 16'd28386, 16'd27984, 16'd43129, 16'd3919}; // indx = 2737
    #10;
    addra = 32'd87616;
    dina = {96'd0, 16'd32388, 16'd17893, 16'd944, 16'd9463, 16'd13555, 16'd28163, 16'd10900, 16'd41562, 16'd16574, 16'd7401}; // indx = 2738
    #10;
    addra = 32'd87648;
    dina = {96'd0, 16'd20056, 16'd33266, 16'd44655, 16'd41326, 16'd8764, 16'd1107, 16'd22096, 16'd32341, 16'd24473, 16'd51217}; // indx = 2739
    #10;
    addra = 32'd87680;
    dina = {96'd0, 16'd8190, 16'd48663, 16'd33718, 16'd46577, 16'd383, 16'd33654, 16'd37664, 16'd43517, 16'd59442, 16'd50828}; // indx = 2740
    #10;
    addra = 32'd87712;
    dina = {96'd0, 16'd26300, 16'd10220, 16'd54785, 16'd5518, 16'd51423, 16'd10001, 16'd19463, 16'd5400, 16'd17511, 16'd25124}; // indx = 2741
    #10;
    addra = 32'd87744;
    dina = {96'd0, 16'd26099, 16'd39259, 16'd42330, 16'd32107, 16'd57777, 16'd38146, 16'd35264, 16'd24318, 16'd46456, 16'd40145}; // indx = 2742
    #10;
    addra = 32'd87776;
    dina = {96'd0, 16'd53462, 16'd55201, 16'd5933, 16'd29894, 16'd19198, 16'd26473, 16'd35111, 16'd53259, 16'd2883, 16'd26695}; // indx = 2743
    #10;
    addra = 32'd87808;
    dina = {96'd0, 16'd695, 16'd59082, 16'd53374, 16'd49410, 16'd30262, 16'd35009, 16'd19141, 16'd21767, 16'd45156, 16'd2271}; // indx = 2744
    #10;
    addra = 32'd87840;
    dina = {96'd0, 16'd7864, 16'd15321, 16'd50715, 16'd35729, 16'd27677, 16'd62756, 16'd33247, 16'd32130, 16'd58774, 16'd1470}; // indx = 2745
    #10;
    addra = 32'd87872;
    dina = {96'd0, 16'd26591, 16'd4027, 16'd46777, 16'd8604, 16'd65487, 16'd1838, 16'd33647, 16'd22639, 16'd18494, 16'd15676}; // indx = 2746
    #10;
    addra = 32'd87904;
    dina = {96'd0, 16'd2744, 16'd50834, 16'd8527, 16'd19260, 16'd52512, 16'd16145, 16'd13977, 16'd41417, 16'd24229, 16'd33579}; // indx = 2747
    #10;
    addra = 32'd87936;
    dina = {96'd0, 16'd56675, 16'd40788, 16'd10674, 16'd3937, 16'd14643, 16'd61714, 16'd23899, 16'd32200, 16'd51936, 16'd5320}; // indx = 2748
    #10;
    addra = 32'd87968;
    dina = {96'd0, 16'd4670, 16'd52409, 16'd63022, 16'd49641, 16'd10192, 16'd62902, 16'd47954, 16'd49629, 16'd53453, 16'd17478}; // indx = 2749
    #10;
    addra = 32'd88000;
    dina = {96'd0, 16'd52440, 16'd21063, 16'd7199, 16'd64060, 16'd55283, 16'd60783, 16'd31185, 16'd46454, 16'd5651, 16'd16263}; // indx = 2750
    #10;
    addra = 32'd88032;
    dina = {96'd0, 16'd64792, 16'd30124, 16'd56392, 16'd33893, 16'd58089, 16'd57712, 16'd57758, 16'd3863, 16'd45651, 16'd54442}; // indx = 2751
    #10;
    addra = 32'd88064;
    dina = {96'd0, 16'd36850, 16'd12339, 16'd31814, 16'd14559, 16'd26160, 16'd10372, 16'd4685, 16'd13914, 16'd9095, 16'd41040}; // indx = 2752
    #10;
    addra = 32'd88096;
    dina = {96'd0, 16'd59383, 16'd33654, 16'd43320, 16'd18422, 16'd21182, 16'd40625, 16'd17543, 16'd31722, 16'd25106, 16'd56533}; // indx = 2753
    #10;
    addra = 32'd88128;
    dina = {96'd0, 16'd29917, 16'd13461, 16'd27012, 16'd44322, 16'd48338, 16'd17315, 16'd22853, 16'd31068, 16'd54585, 16'd9517}; // indx = 2754
    #10;
    addra = 32'd88160;
    dina = {96'd0, 16'd17506, 16'd62038, 16'd17085, 16'd50075, 16'd47368, 16'd41100, 16'd64598, 16'd50144, 16'd35048, 16'd30042}; // indx = 2755
    #10;
    addra = 32'd88192;
    dina = {96'd0, 16'd61049, 16'd529, 16'd41862, 16'd47790, 16'd717, 16'd3203, 16'd5160, 16'd59091, 16'd51407, 16'd3936}; // indx = 2756
    #10;
    addra = 32'd88224;
    dina = {96'd0, 16'd58928, 16'd39124, 16'd56072, 16'd48919, 16'd38881, 16'd15151, 16'd56661, 16'd7045, 16'd57427, 16'd56150}; // indx = 2757
    #10;
    addra = 32'd88256;
    dina = {96'd0, 16'd21469, 16'd19153, 16'd55518, 16'd12551, 16'd64340, 16'd50754, 16'd57904, 16'd58426, 16'd11640, 16'd34259}; // indx = 2758
    #10;
    addra = 32'd88288;
    dina = {96'd0, 16'd36718, 16'd60260, 16'd25832, 16'd29513, 16'd20705, 16'd30792, 16'd64440, 16'd47737, 16'd42589, 16'd16750}; // indx = 2759
    #10;
    addra = 32'd88320;
    dina = {96'd0, 16'd30115, 16'd3719, 16'd26244, 16'd61849, 16'd44128, 16'd39819, 16'd46864, 16'd58834, 16'd35156, 16'd14556}; // indx = 2760
    #10;
    addra = 32'd88352;
    dina = {96'd0, 16'd42814, 16'd30402, 16'd64794, 16'd27406, 16'd1356, 16'd41886, 16'd4180, 16'd20390, 16'd63457, 16'd59768}; // indx = 2761
    #10;
    addra = 32'd88384;
    dina = {96'd0, 16'd23219, 16'd11214, 16'd8019, 16'd30255, 16'd14879, 16'd51601, 16'd4544, 16'd61601, 16'd59362, 16'd64187}; // indx = 2762
    #10;
    addra = 32'd88416;
    dina = {96'd0, 16'd56898, 16'd58752, 16'd13460, 16'd55331, 16'd13205, 16'd64723, 16'd27940, 16'd41611, 16'd64825, 16'd10552}; // indx = 2763
    #10;
    addra = 32'd88448;
    dina = {96'd0, 16'd52705, 16'd52723, 16'd48961, 16'd27817, 16'd25620, 16'd52216, 16'd37594, 16'd61519, 16'd25107, 16'd8356}; // indx = 2764
    #10;
    addra = 32'd88480;
    dina = {96'd0, 16'd23753, 16'd36835, 16'd15812, 16'd29832, 16'd45781, 16'd20633, 16'd40823, 16'd50166, 16'd61421, 16'd49649}; // indx = 2765
    #10;
    addra = 32'd88512;
    dina = {96'd0, 16'd34704, 16'd14718, 16'd25906, 16'd57227, 16'd15192, 16'd2690, 16'd26916, 16'd42221, 16'd8419, 16'd31062}; // indx = 2766
    #10;
    addra = 32'd88544;
    dina = {96'd0, 16'd34425, 16'd8075, 16'd8417, 16'd16176, 16'd4356, 16'd9634, 16'd42942, 16'd13878, 16'd838, 16'd7524}; // indx = 2767
    #10;
    addra = 32'd88576;
    dina = {96'd0, 16'd2408, 16'd50821, 16'd5442, 16'd64876, 16'd17613, 16'd39877, 16'd62573, 16'd30291, 16'd18403, 16'd48738}; // indx = 2768
    #10;
    addra = 32'd88608;
    dina = {96'd0, 16'd19593, 16'd22165, 16'd1471, 16'd6792, 16'd45469, 16'd15488, 16'd43950, 16'd54668, 16'd23338, 16'd1147}; // indx = 2769
    #10;
    addra = 32'd88640;
    dina = {96'd0, 16'd34182, 16'd29103, 16'd24256, 16'd738, 16'd1286, 16'd55671, 16'd29758, 16'd18168, 16'd4830, 16'd14495}; // indx = 2770
    #10;
    addra = 32'd88672;
    dina = {96'd0, 16'd23564, 16'd32814, 16'd11133, 16'd62925, 16'd9101, 16'd54334, 16'd62154, 16'd44168, 16'd612, 16'd17866}; // indx = 2771
    #10;
    addra = 32'd88704;
    dina = {96'd0, 16'd37555, 16'd26440, 16'd64703, 16'd29778, 16'd2418, 16'd48709, 16'd59888, 16'd40796, 16'd4975, 16'd40480}; // indx = 2772
    #10;
    addra = 32'd88736;
    dina = {96'd0, 16'd62967, 16'd15546, 16'd5554, 16'd1360, 16'd3859, 16'd11158, 16'd42494, 16'd48226, 16'd18092, 16'd50630}; // indx = 2773
    #10;
    addra = 32'd88768;
    dina = {96'd0, 16'd35601, 16'd54136, 16'd5479, 16'd1627, 16'd25432, 16'd4414, 16'd38393, 16'd4812, 16'd52475, 16'd57364}; // indx = 2774
    #10;
    addra = 32'd88800;
    dina = {96'd0, 16'd40032, 16'd12518, 16'd6250, 16'd26953, 16'd22522, 16'd51204, 16'd51474, 16'd61510, 16'd40067, 16'd47840}; // indx = 2775
    #10;
    addra = 32'd88832;
    dina = {96'd0, 16'd35786, 16'd59750, 16'd11867, 16'd12991, 16'd16744, 16'd35911, 16'd65258, 16'd45314, 16'd30787, 16'd32698}; // indx = 2776
    #10;
    addra = 32'd88864;
    dina = {96'd0, 16'd41138, 16'd27087, 16'd24373, 16'd25377, 16'd25230, 16'd5272, 16'd23994, 16'd8595, 16'd28960, 16'd28687}; // indx = 2777
    #10;
    addra = 32'd88896;
    dina = {96'd0, 16'd20399, 16'd64458, 16'd52397, 16'd34486, 16'd23467, 16'd9470, 16'd44701, 16'd42666, 16'd24942, 16'd32597}; // indx = 2778
    #10;
    addra = 32'd88928;
    dina = {96'd0, 16'd52441, 16'd48950, 16'd19572, 16'd44936, 16'd25287, 16'd64385, 16'd12210, 16'd1059, 16'd49716, 16'd37085}; // indx = 2779
    #10;
    addra = 32'd88960;
    dina = {96'd0, 16'd59844, 16'd48114, 16'd56194, 16'd25928, 16'd37965, 16'd39130, 16'd37678, 16'd56826, 16'd36637, 16'd51554}; // indx = 2780
    #10;
    addra = 32'd88992;
    dina = {96'd0, 16'd47237, 16'd5903, 16'd53073, 16'd14400, 16'd33024, 16'd55809, 16'd43777, 16'd42808, 16'd51532, 16'd63141}; // indx = 2781
    #10;
    addra = 32'd89024;
    dina = {96'd0, 16'd17815, 16'd19092, 16'd64974, 16'd6512, 16'd27230, 16'd23261, 16'd32089, 16'd10106, 16'd61078, 16'd18023}; // indx = 2782
    #10;
    addra = 32'd89056;
    dina = {96'd0, 16'd64147, 16'd42240, 16'd8977, 16'd11599, 16'd3379, 16'd23517, 16'd41388, 16'd41023, 16'd3221, 16'd41580}; // indx = 2783
    #10;
    addra = 32'd89088;
    dina = {96'd0, 16'd57442, 16'd19124, 16'd2697, 16'd55646, 16'd60668, 16'd22792, 16'd13299, 16'd45495, 16'd29463, 16'd19368}; // indx = 2784
    #10;
    addra = 32'd89120;
    dina = {96'd0, 16'd31211, 16'd38144, 16'd49633, 16'd23686, 16'd8356, 16'd42622, 16'd14163, 16'd48833, 16'd37530, 16'd936}; // indx = 2785
    #10;
    addra = 32'd89152;
    dina = {96'd0, 16'd32986, 16'd11654, 16'd32851, 16'd42127, 16'd58182, 16'd25523, 16'd24689, 16'd43781, 16'd41137, 16'd61876}; // indx = 2786
    #10;
    addra = 32'd89184;
    dina = {96'd0, 16'd64981, 16'd8590, 16'd31562, 16'd47224, 16'd48881, 16'd49365, 16'd5909, 16'd48778, 16'd31378, 16'd43435}; // indx = 2787
    #10;
    addra = 32'd89216;
    dina = {96'd0, 16'd47605, 16'd23744, 16'd53618, 16'd32968, 16'd327, 16'd44400, 16'd5567, 16'd1064, 16'd37378, 16'd17847}; // indx = 2788
    #10;
    addra = 32'd89248;
    dina = {96'd0, 16'd52239, 16'd46640, 16'd34116, 16'd3879, 16'd40190, 16'd7306, 16'd49157, 16'd31827, 16'd51820, 16'd45889}; // indx = 2789
    #10;
    addra = 32'd89280;
    dina = {96'd0, 16'd48392, 16'd26392, 16'd33095, 16'd20642, 16'd56273, 16'd4025, 16'd27653, 16'd48193, 16'd53198, 16'd30716}; // indx = 2790
    #10;
    addra = 32'd89312;
    dina = {96'd0, 16'd5318, 16'd34947, 16'd45412, 16'd43434, 16'd5737, 16'd28402, 16'd23547, 16'd54974, 16'd28489, 16'd11311}; // indx = 2791
    #10;
    addra = 32'd89344;
    dina = {96'd0, 16'd42293, 16'd50853, 16'd9488, 16'd47054, 16'd7, 16'd11382, 16'd51498, 16'd42628, 16'd35059, 16'd31823}; // indx = 2792
    #10;
    addra = 32'd89376;
    dina = {96'd0, 16'd3998, 16'd13769, 16'd51599, 16'd59786, 16'd50065, 16'd61596, 16'd44905, 16'd35459, 16'd45551, 16'd59164}; // indx = 2793
    #10;
    addra = 32'd89408;
    dina = {96'd0, 16'd14491, 16'd17068, 16'd23134, 16'd17825, 16'd41163, 16'd27247, 16'd62797, 16'd49226, 16'd63252, 16'd10988}; // indx = 2794
    #10;
    addra = 32'd89440;
    dina = {96'd0, 16'd39688, 16'd11352, 16'd22565, 16'd2089, 16'd8557, 16'd28519, 16'd18424, 16'd49832, 16'd57041, 16'd56699}; // indx = 2795
    #10;
    addra = 32'd89472;
    dina = {96'd0, 16'd33264, 16'd3581, 16'd56017, 16'd12767, 16'd47219, 16'd63009, 16'd5324, 16'd22982, 16'd29521, 16'd12129}; // indx = 2796
    #10;
    addra = 32'd89504;
    dina = {96'd0, 16'd54028, 16'd40141, 16'd29884, 16'd42789, 16'd28335, 16'd43038, 16'd57756, 16'd30083, 16'd42060, 16'd24332}; // indx = 2797
    #10;
    addra = 32'd89536;
    dina = {96'd0, 16'd27137, 16'd14629, 16'd4916, 16'd56314, 16'd35107, 16'd46889, 16'd3462, 16'd16349, 16'd49696, 16'd23619}; // indx = 2798
    #10;
    addra = 32'd89568;
    dina = {96'd0, 16'd46006, 16'd39019, 16'd27799, 16'd13472, 16'd16680, 16'd10979, 16'd20043, 16'd63042, 16'd30960, 16'd53299}; // indx = 2799
    #10;
    addra = 32'd89600;
    dina = {96'd0, 16'd38446, 16'd9501, 16'd4349, 16'd55224, 16'd4001, 16'd31136, 16'd58015, 16'd3157, 16'd47701, 16'd23481}; // indx = 2800
    #10;
    addra = 32'd89632;
    dina = {96'd0, 16'd17956, 16'd52660, 16'd35716, 16'd8639, 16'd8612, 16'd63804, 16'd42685, 16'd30004, 16'd27624, 16'd8973}; // indx = 2801
    #10;
    addra = 32'd89664;
    dina = {96'd0, 16'd50090, 16'd27658, 16'd58388, 16'd39878, 16'd61086, 16'd34679, 16'd50147, 16'd568, 16'd40027, 16'd55647}; // indx = 2802
    #10;
    addra = 32'd89696;
    dina = {96'd0, 16'd55317, 16'd46118, 16'd15600, 16'd65182, 16'd44478, 16'd24548, 16'd12237, 16'd540, 16'd57781, 16'd44977}; // indx = 2803
    #10;
    addra = 32'd89728;
    dina = {96'd0, 16'd31149, 16'd514, 16'd14691, 16'd54717, 16'd15487, 16'd54123, 16'd40497, 16'd40416, 16'd56078, 16'd28473}; // indx = 2804
    #10;
    addra = 32'd89760;
    dina = {96'd0, 16'd15842, 16'd43582, 16'd51958, 16'd62237, 16'd2550, 16'd30441, 16'd50302, 16'd34406, 16'd24974, 16'd20888}; // indx = 2805
    #10;
    addra = 32'd89792;
    dina = {96'd0, 16'd22079, 16'd29732, 16'd65091, 16'd44691, 16'd13784, 16'd23244, 16'd10000, 16'd48441, 16'd9203, 16'd54625}; // indx = 2806
    #10;
    addra = 32'd89824;
    dina = {96'd0, 16'd24961, 16'd35140, 16'd1085, 16'd16548, 16'd37141, 16'd36254, 16'd55171, 16'd18432, 16'd10966, 16'd18260}; // indx = 2807
    #10;
    addra = 32'd89856;
    dina = {96'd0, 16'd53199, 16'd37824, 16'd50501, 16'd11434, 16'd30013, 16'd37266, 16'd28386, 16'd9109, 16'd44308, 16'd7087}; // indx = 2808
    #10;
    addra = 32'd89888;
    dina = {96'd0, 16'd53348, 16'd39993, 16'd8461, 16'd30973, 16'd55887, 16'd16057, 16'd22858, 16'd21568, 16'd43917, 16'd59193}; // indx = 2809
    #10;
    addra = 32'd89920;
    dina = {96'd0, 16'd9144, 16'd6497, 16'd42997, 16'd2368, 16'd64921, 16'd13836, 16'd13823, 16'd7459, 16'd29848, 16'd39558}; // indx = 2810
    #10;
    addra = 32'd89952;
    dina = {96'd0, 16'd40095, 16'd2157, 16'd6055, 16'd53601, 16'd3238, 16'd26441, 16'd44518, 16'd27243, 16'd24799, 16'd2398}; // indx = 2811
    #10;
    addra = 32'd89984;
    dina = {96'd0, 16'd57522, 16'd51113, 16'd29177, 16'd31149, 16'd31343, 16'd13740, 16'd52417, 16'd17772, 16'd58230, 16'd6551}; // indx = 2812
    #10;
    addra = 32'd90016;
    dina = {96'd0, 16'd3618, 16'd15986, 16'd52017, 16'd35862, 16'd33583, 16'd41619, 16'd38634, 16'd49436, 16'd38033, 16'd28101}; // indx = 2813
    #10;
    addra = 32'd90048;
    dina = {96'd0, 16'd20182, 16'd61087, 16'd32647, 16'd7424, 16'd32626, 16'd51024, 16'd14282, 16'd64563, 16'd60247, 16'd1206}; // indx = 2814
    #10;
    addra = 32'd90080;
    dina = {96'd0, 16'd34181, 16'd33742, 16'd3950, 16'd50713, 16'd53281, 16'd25433, 16'd43293, 16'd19469, 16'd54978, 16'd38307}; // indx = 2815
    #10;
    addra = 32'd90112;
    dina = {96'd0, 16'd32062, 16'd3798, 16'd41866, 16'd40964, 16'd58240, 16'd38672, 16'd28495, 16'd64913, 16'd47568, 16'd452}; // indx = 2816
    #10;
    addra = 32'd90144;
    dina = {96'd0, 16'd12237, 16'd46976, 16'd59321, 16'd19918, 16'd30697, 16'd25642, 16'd41124, 16'd34467, 16'd21936, 16'd6766}; // indx = 2817
    #10;
    addra = 32'd90176;
    dina = {96'd0, 16'd13787, 16'd8598, 16'd64906, 16'd19580, 16'd26084, 16'd55943, 16'd11975, 16'd37660, 16'd63059, 16'd62825}; // indx = 2818
    #10;
    addra = 32'd90208;
    dina = {96'd0, 16'd2746, 16'd3573, 16'd17306, 16'd20617, 16'd62851, 16'd50469, 16'd26105, 16'd39383, 16'd21466, 16'd62285}; // indx = 2819
    #10;
    addra = 32'd90240;
    dina = {96'd0, 16'd31776, 16'd14491, 16'd13057, 16'd19841, 16'd59100, 16'd15417, 16'd61420, 16'd34200, 16'd48299, 16'd30364}; // indx = 2820
    #10;
    addra = 32'd90272;
    dina = {96'd0, 16'd52620, 16'd15312, 16'd38577, 16'd2188, 16'd45249, 16'd51266, 16'd35339, 16'd59110, 16'd54767, 16'd27970}; // indx = 2821
    #10;
    addra = 32'd90304;
    dina = {96'd0, 16'd7328, 16'd55339, 16'd61168, 16'd52382, 16'd31637, 16'd31391, 16'd9600, 16'd16185, 16'd1987, 16'd42502}; // indx = 2822
    #10;
    addra = 32'd90336;
    dina = {96'd0, 16'd58571, 16'd4872, 16'd24865, 16'd58432, 16'd25036, 16'd9048, 16'd6434, 16'd59025, 16'd1831, 16'd34888}; // indx = 2823
    #10;
    addra = 32'd90368;
    dina = {96'd0, 16'd4375, 16'd9653, 16'd60667, 16'd5018, 16'd59192, 16'd1437, 16'd62264, 16'd59562, 16'd15770, 16'd17255}; // indx = 2824
    #10;
    addra = 32'd90400;
    dina = {96'd0, 16'd9569, 16'd22376, 16'd40733, 16'd28605, 16'd42358, 16'd20406, 16'd21767, 16'd35993, 16'd33044, 16'd13030}; // indx = 2825
    #10;
    addra = 32'd90432;
    dina = {96'd0, 16'd30212, 16'd60895, 16'd16100, 16'd11238, 16'd54658, 16'd20689, 16'd15418, 16'd55148, 16'd28748, 16'd6738}; // indx = 2826
    #10;
    addra = 32'd90464;
    dina = {96'd0, 16'd26773, 16'd5665, 16'd41759, 16'd61591, 16'd34062, 16'd27342, 16'd60021, 16'd35264, 16'd33276, 16'd56708}; // indx = 2827
    #10;
    addra = 32'd90496;
    dina = {96'd0, 16'd27851, 16'd16137, 16'd12272, 16'd31252, 16'd24182, 16'd6658, 16'd17129, 16'd61682, 16'd3982, 16'd15644}; // indx = 2828
    #10;
    addra = 32'd90528;
    dina = {96'd0, 16'd27513, 16'd44999, 16'd10210, 16'd15234, 16'd45951, 16'd52798, 16'd45921, 16'd35364, 16'd63996, 16'd58767}; // indx = 2829
    #10;
    addra = 32'd90560;
    dina = {96'd0, 16'd30863, 16'd17799, 16'd9572, 16'd59461, 16'd8282, 16'd62584, 16'd50777, 16'd56018, 16'd53531, 16'd7920}; // indx = 2830
    #10;
    addra = 32'd90592;
    dina = {96'd0, 16'd24133, 16'd16089, 16'd15387, 16'd57744, 16'd56977, 16'd50345, 16'd39466, 16'd12686, 16'd49570, 16'd55129}; // indx = 2831
    #10;
    addra = 32'd90624;
    dina = {96'd0, 16'd64573, 16'd60638, 16'd21015, 16'd48118, 16'd47549, 16'd33396, 16'd3584, 16'd39700, 16'd6895, 16'd30292}; // indx = 2832
    #10;
    addra = 32'd90656;
    dina = {96'd0, 16'd33588, 16'd14894, 16'd22085, 16'd45527, 16'd29216, 16'd5474, 16'd63492, 16'd3035, 16'd4713, 16'd21010}; // indx = 2833
    #10;
    addra = 32'd90688;
    dina = {96'd0, 16'd27266, 16'd54145, 16'd16873, 16'd17317, 16'd80, 16'd58818, 16'd3405, 16'd20404, 16'd35031, 16'd61479}; // indx = 2834
    #10;
    addra = 32'd90720;
    dina = {96'd0, 16'd60270, 16'd59879, 16'd34746, 16'd46989, 16'd49950, 16'd28167, 16'd3827, 16'd41744, 16'd23508, 16'd30693}; // indx = 2835
    #10;
    addra = 32'd90752;
    dina = {96'd0, 16'd42830, 16'd29344, 16'd855, 16'd58468, 16'd51702, 16'd29828, 16'd21108, 16'd32599, 16'd40402, 16'd48486}; // indx = 2836
    #10;
    addra = 32'd90784;
    dina = {96'd0, 16'd53969, 16'd46571, 16'd31187, 16'd14869, 16'd58237, 16'd46288, 16'd923, 16'd48439, 16'd55810, 16'd4218}; // indx = 2837
    #10;
    addra = 32'd90816;
    dina = {96'd0, 16'd7749, 16'd58511, 16'd27615, 16'd49993, 16'd33111, 16'd4320, 16'd65470, 16'd41399, 16'd42049, 16'd30629}; // indx = 2838
    #10;
    addra = 32'd90848;
    dina = {96'd0, 16'd57422, 16'd22292, 16'd28630, 16'd1294, 16'd9171, 16'd45928, 16'd23581, 16'd35661, 16'd63729, 16'd27773}; // indx = 2839
    #10;
    addra = 32'd90880;
    dina = {96'd0, 16'd21833, 16'd18438, 16'd17782, 16'd6081, 16'd32581, 16'd45750, 16'd13782, 16'd27302, 16'd9622, 16'd6132}; // indx = 2840
    #10;
    addra = 32'd90912;
    dina = {96'd0, 16'd62994, 16'd53472, 16'd10550, 16'd13748, 16'd56719, 16'd5523, 16'd53576, 16'd59107, 16'd29580, 16'd22678}; // indx = 2841
    #10;
    addra = 32'd90944;
    dina = {96'd0, 16'd62180, 16'd54423, 16'd11701, 16'd26038, 16'd16099, 16'd41415, 16'd41485, 16'd61984, 16'd62134, 16'd28316}; // indx = 2842
    #10;
    addra = 32'd90976;
    dina = {96'd0, 16'd9973, 16'd60570, 16'd12886, 16'd37644, 16'd58398, 16'd37235, 16'd12190, 16'd34779, 16'd30203, 16'd59126}; // indx = 2843
    #10;
    addra = 32'd91008;
    dina = {96'd0, 16'd19471, 16'd22455, 16'd63783, 16'd41591, 16'd54307, 16'd11503, 16'd57498, 16'd62084, 16'd53096, 16'd25899}; // indx = 2844
    #10;
    addra = 32'd91040;
    dina = {96'd0, 16'd31018, 16'd60781, 16'd61613, 16'd18072, 16'd29127, 16'd25090, 16'd21804, 16'd22369, 16'd16059, 16'd63462}; // indx = 2845
    #10;
    addra = 32'd91072;
    dina = {96'd0, 16'd204, 16'd37606, 16'd46196, 16'd35107, 16'd10288, 16'd23105, 16'd35540, 16'd1393, 16'd47799, 16'd64627}; // indx = 2846
    #10;
    addra = 32'd91104;
    dina = {96'd0, 16'd51696, 16'd38473, 16'd39708, 16'd32643, 16'd14072, 16'd51997, 16'd30631, 16'd44632, 16'd32342, 16'd17635}; // indx = 2847
    #10;
    addra = 32'd91136;
    dina = {96'd0, 16'd29332, 16'd17640, 16'd7856, 16'd40545, 16'd29490, 16'd19450, 16'd37428, 16'd29726, 16'd20923, 16'd12365}; // indx = 2848
    #10;
    addra = 32'd91168;
    dina = {96'd0, 16'd56610, 16'd42746, 16'd63152, 16'd6437, 16'd34200, 16'd14605, 16'd2555, 16'd49836, 16'd23774, 16'd42366}; // indx = 2849
    #10;
    addra = 32'd91200;
    dina = {96'd0, 16'd55347, 16'd20901, 16'd25148, 16'd59662, 16'd19334, 16'd52897, 16'd62473, 16'd58, 16'd3906, 16'd27008}; // indx = 2850
    #10;
    addra = 32'd91232;
    dina = {96'd0, 16'd35602, 16'd4685, 16'd50210, 16'd57687, 16'd56193, 16'd47325, 16'd38961, 16'd49476, 16'd64424, 16'd150}; // indx = 2851
    #10;
    addra = 32'd91264;
    dina = {96'd0, 16'd65040, 16'd54204, 16'd23735, 16'd43787, 16'd41824, 16'd36075, 16'd43923, 16'd64293, 16'd65318, 16'd5785}; // indx = 2852
    #10;
    addra = 32'd91296;
    dina = {96'd0, 16'd27053, 16'd59229, 16'd39693, 16'd24844, 16'd27668, 16'd64977, 16'd16336, 16'd25818, 16'd43871, 16'd41895}; // indx = 2853
    #10;
    addra = 32'd91328;
    dina = {96'd0, 16'd20874, 16'd1072, 16'd46322, 16'd54363, 16'd28474, 16'd28682, 16'd49625, 16'd18111, 16'd32250, 16'd38838}; // indx = 2854
    #10;
    addra = 32'd91360;
    dina = {96'd0, 16'd59128, 16'd64785, 16'd64772, 16'd49448, 16'd20806, 16'd8822, 16'd1437, 16'd27419, 16'd48197, 16'd17894}; // indx = 2855
    #10;
    addra = 32'd91392;
    dina = {96'd0, 16'd39056, 16'd35585, 16'd61060, 16'd41873, 16'd26363, 16'd55369, 16'd64661, 16'd40000, 16'd21539, 16'd3411}; // indx = 2856
    #10;
    addra = 32'd91424;
    dina = {96'd0, 16'd58760, 16'd47500, 16'd55829, 16'd40956, 16'd54556, 16'd53755, 16'd50041, 16'd7389, 16'd32749, 16'd64855}; // indx = 2857
    #10;
    addra = 32'd91456;
    dina = {96'd0, 16'd34496, 16'd53577, 16'd51002, 16'd12624, 16'd42595, 16'd40037, 16'd15327, 16'd11197, 16'd63882, 16'd27116}; // indx = 2858
    #10;
    addra = 32'd91488;
    dina = {96'd0, 16'd16882, 16'd17075, 16'd30667, 16'd35685, 16'd41887, 16'd56581, 16'd3739, 16'd15426, 16'd62652, 16'd60433}; // indx = 2859
    #10;
    addra = 32'd91520;
    dina = {96'd0, 16'd64252, 16'd61378, 16'd50737, 16'd29593, 16'd42549, 16'd49938, 16'd40295, 16'd17936, 16'd40267, 16'd35011}; // indx = 2860
    #10;
    addra = 32'd91552;
    dina = {96'd0, 16'd53109, 16'd18198, 16'd27350, 16'd49511, 16'd24796, 16'd18124, 16'd60259, 16'd17514, 16'd51795, 16'd39561}; // indx = 2861
    #10;
    addra = 32'd91584;
    dina = {96'd0, 16'd58401, 16'd25731, 16'd46600, 16'd55490, 16'd23450, 16'd23616, 16'd39344, 16'd20298, 16'd48588, 16'd45290}; // indx = 2862
    #10;
    addra = 32'd91616;
    dina = {96'd0, 16'd54105, 16'd17173, 16'd58454, 16'd60277, 16'd52282, 16'd40347, 16'd42938, 16'd16494, 16'd57513, 16'd15608}; // indx = 2863
    #10;
    addra = 32'd91648;
    dina = {96'd0, 16'd59416, 16'd28762, 16'd8170, 16'd64647, 16'd29762, 16'd13721, 16'd59237, 16'd63257, 16'd5724, 16'd46625}; // indx = 2864
    #10;
    addra = 32'd91680;
    dina = {96'd0, 16'd55331, 16'd19900, 16'd57524, 16'd46455, 16'd35948, 16'd19737, 16'd43119, 16'd60062, 16'd54369, 16'd47052}; // indx = 2865
    #10;
    addra = 32'd91712;
    dina = {96'd0, 16'd40158, 16'd9264, 16'd11310, 16'd50038, 16'd36363, 16'd28846, 16'd9155, 16'd35304, 16'd50710, 16'd45231}; // indx = 2866
    #10;
    addra = 32'd91744;
    dina = {96'd0, 16'd17695, 16'd29527, 16'd10315, 16'd12048, 16'd61873, 16'd33196, 16'd31683, 16'd14829, 16'd9402, 16'd45900}; // indx = 2867
    #10;
    addra = 32'd91776;
    dina = {96'd0, 16'd33014, 16'd22449, 16'd27009, 16'd40894, 16'd52326, 16'd14967, 16'd51521, 16'd17810, 16'd6793, 16'd32473}; // indx = 2868
    #10;
    addra = 32'd91808;
    dina = {96'd0, 16'd19698, 16'd48711, 16'd31251, 16'd17973, 16'd54454, 16'd26737, 16'd19968, 16'd5314, 16'd3453, 16'd35952}; // indx = 2869
    #10;
    addra = 32'd91840;
    dina = {96'd0, 16'd32059, 16'd39628, 16'd45791, 16'd9858, 16'd28730, 16'd26022, 16'd35348, 16'd1715, 16'd1592, 16'd16505}; // indx = 2870
    #10;
    addra = 32'd91872;
    dina = {96'd0, 16'd57656, 16'd19030, 16'd52526, 16'd13613, 16'd44527, 16'd35000, 16'd45019, 16'd30963, 16'd43711, 16'd57171}; // indx = 2871
    #10;
    addra = 32'd91904;
    dina = {96'd0, 16'd11676, 16'd42547, 16'd45665, 16'd21518, 16'd43918, 16'd7793, 16'd52630, 16'd54531, 16'd58079, 16'd11233}; // indx = 2872
    #10;
    addra = 32'd91936;
    dina = {96'd0, 16'd44373, 16'd46621, 16'd9257, 16'd28207, 16'd49332, 16'd39230, 16'd4835, 16'd19511, 16'd48836, 16'd19605}; // indx = 2873
    #10;
    addra = 32'd91968;
    dina = {96'd0, 16'd24505, 16'd0, 16'd28094, 16'd49691, 16'd53436, 16'd40962, 16'd58464, 16'd17955, 16'd26482, 16'd59756}; // indx = 2874
    #10;
    addra = 32'd92000;
    dina = {96'd0, 16'd28185, 16'd23718, 16'd7370, 16'd41619, 16'd64918, 16'd53401, 16'd48684, 16'd46752, 16'd11614, 16'd46023}; // indx = 2875
    #10;
    addra = 32'd92032;
    dina = {96'd0, 16'd50760, 16'd45455, 16'd64930, 16'd10403, 16'd590, 16'd63409, 16'd16098, 16'd46716, 16'd46459, 16'd54765}; // indx = 2876
    #10;
    addra = 32'd92064;
    dina = {96'd0, 16'd36609, 16'd23760, 16'd59792, 16'd25099, 16'd11115, 16'd13225, 16'd45574, 16'd56308, 16'd33495, 16'd45038}; // indx = 2877
    #10;
    addra = 32'd92096;
    dina = {96'd0, 16'd50503, 16'd22162, 16'd47545, 16'd22065, 16'd34711, 16'd55422, 16'd9529, 16'd4081, 16'd2565, 16'd6191}; // indx = 2878
    #10;
    addra = 32'd92128;
    dina = {96'd0, 16'd23568, 16'd62011, 16'd4765, 16'd64247, 16'd34895, 16'd62615, 16'd23763, 16'd20794, 16'd60473, 16'd2596}; // indx = 2879
    #10;
    addra = 32'd92160;
    dina = {96'd0, 16'd3481, 16'd18071, 16'd1911, 16'd49190, 16'd5126, 16'd23082, 16'd40056, 16'd60451, 16'd23714, 16'd33244}; // indx = 2880
    #10;
    addra = 32'd92192;
    dina = {96'd0, 16'd39167, 16'd63223, 16'd49386, 16'd54729, 16'd14548, 16'd51313, 16'd52609, 16'd32955, 16'd38862, 16'd39612}; // indx = 2881
    #10;
    addra = 32'd92224;
    dina = {96'd0, 16'd20303, 16'd63441, 16'd62010, 16'd3107, 16'd28831, 16'd30165, 16'd6853, 16'd36110, 16'd50236, 16'd18199}; // indx = 2882
    #10;
    addra = 32'd92256;
    dina = {96'd0, 16'd24311, 16'd13225, 16'd16870, 16'd34468, 16'd10112, 16'd41576, 16'd31505, 16'd20905, 16'd62663, 16'd34000}; // indx = 2883
    #10;
    addra = 32'd92288;
    dina = {96'd0, 16'd19388, 16'd29460, 16'd61773, 16'd27312, 16'd58477, 16'd55456, 16'd3903, 16'd52116, 16'd64474, 16'd510}; // indx = 2884
    #10;
    addra = 32'd92320;
    dina = {96'd0, 16'd23230, 16'd15010, 16'd2250, 16'd51663, 16'd30449, 16'd63792, 16'd15298, 16'd27734, 16'd15620, 16'd50188}; // indx = 2885
    #10;
    addra = 32'd92352;
    dina = {96'd0, 16'd11630, 16'd34288, 16'd41157, 16'd15790, 16'd17248, 16'd31672, 16'd22978, 16'd22100, 16'd35114, 16'd15505}; // indx = 2886
    #10;
    addra = 32'd92384;
    dina = {96'd0, 16'd30796, 16'd57101, 16'd27714, 16'd43068, 16'd62555, 16'd60405, 16'd9037, 16'd23464, 16'd55743, 16'd19348}; // indx = 2887
    #10;
    addra = 32'd92416;
    dina = {96'd0, 16'd7087, 16'd6093, 16'd62934, 16'd9249, 16'd62274, 16'd32739, 16'd52992, 16'd29863, 16'd10360, 16'd29264}; // indx = 2888
    #10;
    addra = 32'd92448;
    dina = {96'd0, 16'd33209, 16'd61404, 16'd56957, 16'd16311, 16'd13259, 16'd234, 16'd805, 16'd57452, 16'd62448, 16'd4682}; // indx = 2889
    #10;
    addra = 32'd92480;
    dina = {96'd0, 16'd23905, 16'd19135, 16'd51927, 16'd3392, 16'd60766, 16'd8114, 16'd22410, 16'd4981, 16'd445, 16'd51240}; // indx = 2890
    #10;
    addra = 32'd92512;
    dina = {96'd0, 16'd709, 16'd56254, 16'd6079, 16'd54239, 16'd18162, 16'd60420, 16'd6543, 16'd11372, 16'd6288, 16'd33809}; // indx = 2891
    #10;
    addra = 32'd92544;
    dina = {96'd0, 16'd64905, 16'd22364, 16'd27914, 16'd47732, 16'd29818, 16'd19826, 16'd21002, 16'd16471, 16'd53630, 16'd7115}; // indx = 2892
    #10;
    addra = 32'd92576;
    dina = {96'd0, 16'd8965, 16'd52546, 16'd64334, 16'd46258, 16'd5772, 16'd33635, 16'd20206, 16'd2770, 16'd9692, 16'd38187}; // indx = 2893
    #10;
    addra = 32'd92608;
    dina = {96'd0, 16'd28048, 16'd37994, 16'd48859, 16'd27169, 16'd32467, 16'd64655, 16'd35300, 16'd1438, 16'd64710, 16'd7707}; // indx = 2894
    #10;
    addra = 32'd92640;
    dina = {96'd0, 16'd19292, 16'd8787, 16'd29820, 16'd35611, 16'd15974, 16'd9, 16'd24943, 16'd5936, 16'd13708, 16'd43659}; // indx = 2895
    #10;
    addra = 32'd92672;
    dina = {96'd0, 16'd41451, 16'd4095, 16'd24097, 16'd19225, 16'd60863, 16'd23165, 16'd55803, 16'd20056, 16'd48515, 16'd59955}; // indx = 2896
    #10;
    addra = 32'd92704;
    dina = {96'd0, 16'd27153, 16'd55337, 16'd25276, 16'd62641, 16'd5279, 16'd43539, 16'd21543, 16'd9307, 16'd28600, 16'd59697}; // indx = 2897
    #10;
    addra = 32'd92736;
    dina = {96'd0, 16'd32629, 16'd2077, 16'd61464, 16'd9696, 16'd2017, 16'd8440, 16'd47672, 16'd62136, 16'd22638, 16'd38582}; // indx = 2898
    #10;
    addra = 32'd92768;
    dina = {96'd0, 16'd19016, 16'd28342, 16'd1806, 16'd6990, 16'd13883, 16'd19037, 16'd2508, 16'd54822, 16'd19880, 16'd2108}; // indx = 2899
    #10;
    addra = 32'd92800;
    dina = {96'd0, 16'd33994, 16'd64652, 16'd24458, 16'd27606, 16'd27043, 16'd5065, 16'd44623, 16'd21248, 16'd10902, 16'd28325}; // indx = 2900
    #10;
    addra = 32'd92832;
    dina = {96'd0, 16'd45381, 16'd35740, 16'd43011, 16'd33140, 16'd3697, 16'd57737, 16'd61021, 16'd29412, 16'd59917, 16'd52839}; // indx = 2901
    #10;
    addra = 32'd92864;
    dina = {96'd0, 16'd22289, 16'd26319, 16'd34739, 16'd18739, 16'd43917, 16'd56137, 16'd51971, 16'd37269, 16'd54681, 16'd6435}; // indx = 2902
    #10;
    addra = 32'd92896;
    dina = {96'd0, 16'd63840, 16'd14195, 16'd39713, 16'd11250, 16'd6430, 16'd53285, 16'd35533, 16'd64123, 16'd37412, 16'd63422}; // indx = 2903
    #10;
    addra = 32'd92928;
    dina = {96'd0, 16'd53585, 16'd44455, 16'd20885, 16'd7136, 16'd49465, 16'd40937, 16'd14801, 16'd4033, 16'd23748, 16'd37206}; // indx = 2904
    #10;
    addra = 32'd92960;
    dina = {96'd0, 16'd42014, 16'd62048, 16'd36384, 16'd50937, 16'd43665, 16'd44059, 16'd12847, 16'd33148, 16'd64185, 16'd37468}; // indx = 2905
    #10;
    addra = 32'd92992;
    dina = {96'd0, 16'd59797, 16'd12539, 16'd14684, 16'd26784, 16'd19258, 16'd21714, 16'd3759, 16'd62247, 16'd1386, 16'd64290}; // indx = 2906
    #10;
    addra = 32'd93024;
    dina = {96'd0, 16'd299, 16'd10318, 16'd14474, 16'd27137, 16'd23718, 16'd39573, 16'd37323, 16'd10086, 16'd44809, 16'd42776}; // indx = 2907
    #10;
    addra = 32'd93056;
    dina = {96'd0, 16'd64533, 16'd6029, 16'd46364, 16'd23568, 16'd60255, 16'd54346, 16'd17413, 16'd15525, 16'd33103, 16'd51873}; // indx = 2908
    #10;
    addra = 32'd93088;
    dina = {96'd0, 16'd48940, 16'd55837, 16'd29358, 16'd23207, 16'd62980, 16'd44223, 16'd42543, 16'd9818, 16'd6751, 16'd12686}; // indx = 2909
    #10;
    addra = 32'd93120;
    dina = {96'd0, 16'd59786, 16'd15096, 16'd46320, 16'd26134, 16'd61109, 16'd35474, 16'd63074, 16'd22356, 16'd9606, 16'd56731}; // indx = 2910
    #10;
    addra = 32'd93152;
    dina = {96'd0, 16'd31633, 16'd35773, 16'd25380, 16'd23782, 16'd4024, 16'd10932, 16'd19681, 16'd22675, 16'd53616, 16'd26484}; // indx = 2911
    #10;
    addra = 32'd93184;
    dina = {96'd0, 16'd41564, 16'd24414, 16'd60189, 16'd8974, 16'd47062, 16'd16080, 16'd17454, 16'd16095, 16'd54837, 16'd27578}; // indx = 2912
    #10;
    addra = 32'd93216;
    dina = {96'd0, 16'd9139, 16'd54331, 16'd3378, 16'd30676, 16'd14003, 16'd30395, 16'd14019, 16'd26526, 16'd32812, 16'd33015}; // indx = 2913
    #10;
    addra = 32'd93248;
    dina = {96'd0, 16'd18588, 16'd59995, 16'd10254, 16'd18594, 16'd19419, 16'd6853, 16'd54465, 16'd17408, 16'd18701, 16'd3740}; // indx = 2914
    #10;
    addra = 32'd93280;
    dina = {96'd0, 16'd43551, 16'd51333, 16'd35075, 16'd25638, 16'd22726, 16'd2099, 16'd22238, 16'd28524, 16'd64268, 16'd65231}; // indx = 2915
    #10;
    addra = 32'd93312;
    dina = {96'd0, 16'd56771, 16'd58872, 16'd35936, 16'd52822, 16'd30520, 16'd65120, 16'd12979, 16'd44696, 16'd16709, 16'd21704}; // indx = 2916
    #10;
    addra = 32'd93344;
    dina = {96'd0, 16'd4995, 16'd14551, 16'd38951, 16'd21355, 16'd19642, 16'd50272, 16'd57393, 16'd16862, 16'd60184, 16'd41983}; // indx = 2917
    #10;
    addra = 32'd93376;
    dina = {96'd0, 16'd32822, 16'd55618, 16'd8325, 16'd588, 16'd50263, 16'd24381, 16'd16042, 16'd30163, 16'd11863, 16'd28846}; // indx = 2918
    #10;
    addra = 32'd93408;
    dina = {96'd0, 16'd55248, 16'd56924, 16'd44105, 16'd62058, 16'd31600, 16'd58184, 16'd12996, 16'd34340, 16'd22269, 16'd24515}; // indx = 2919
    #10;
    addra = 32'd93440;
    dina = {96'd0, 16'd53038, 16'd12520, 16'd60756, 16'd5271, 16'd61054, 16'd45363, 16'd21471, 16'd20164, 16'd22779, 16'd38439}; // indx = 2920
    #10;
    addra = 32'd93472;
    dina = {96'd0, 16'd24360, 16'd64862, 16'd3626, 16'd26297, 16'd33958, 16'd21504, 16'd64720, 16'd20677, 16'd28761, 16'd16266}; // indx = 2921
    #10;
    addra = 32'd93504;
    dina = {96'd0, 16'd45965, 16'd31593, 16'd7673, 16'd65035, 16'd28862, 16'd32600, 16'd2984, 16'd7498, 16'd29217, 16'd22874}; // indx = 2922
    #10;
    addra = 32'd93536;
    dina = {96'd0, 16'd34665, 16'd56014, 16'd55888, 16'd15612, 16'd54025, 16'd64036, 16'd45836, 16'd37477, 16'd57540, 16'd40437}; // indx = 2923
    #10;
    addra = 32'd93568;
    dina = {96'd0, 16'd41493, 16'd48497, 16'd51875, 16'd56051, 16'd7542, 16'd34133, 16'd65008, 16'd15047, 16'd60232, 16'd19846}; // indx = 2924
    #10;
    addra = 32'd93600;
    dina = {96'd0, 16'd56163, 16'd28169, 16'd47219, 16'd27877, 16'd24718, 16'd31871, 16'd21728, 16'd50759, 16'd41500, 16'd51351}; // indx = 2925
    #10;
    addra = 32'd93632;
    dina = {96'd0, 16'd15278, 16'd50653, 16'd264, 16'd58471, 16'd44614, 16'd30262, 16'd52491, 16'd30419, 16'd26820, 16'd57075}; // indx = 2926
    #10;
    addra = 32'd93664;
    dina = {96'd0, 16'd55168, 16'd15236, 16'd59890, 16'd3099, 16'd28023, 16'd19553, 16'd54245, 16'd7741, 16'd57228, 16'd29017}; // indx = 2927
    #10;
    addra = 32'd93696;
    dina = {96'd0, 16'd48971, 16'd64487, 16'd35145, 16'd62991, 16'd45996, 16'd25859, 16'd51225, 16'd55321, 16'd55497, 16'd65179}; // indx = 2928
    #10;
    addra = 32'd93728;
    dina = {96'd0, 16'd24308, 16'd64487, 16'd50887, 16'd20275, 16'd56566, 16'd39482, 16'd42759, 16'd23317, 16'd45200, 16'd6395}; // indx = 2929
    #10;
    addra = 32'd93760;
    dina = {96'd0, 16'd13543, 16'd56900, 16'd55622, 16'd20091, 16'd58159, 16'd41913, 16'd28502, 16'd64644, 16'd50895, 16'd40343}; // indx = 2930
    #10;
    addra = 32'd93792;
    dina = {96'd0, 16'd44019, 16'd56593, 16'd27862, 16'd6449, 16'd46469, 16'd64891, 16'd46181, 16'd53887, 16'd60422, 16'd39357}; // indx = 2931
    #10;
    addra = 32'd93824;
    dina = {96'd0, 16'd8845, 16'd3118, 16'd1170, 16'd10977, 16'd63399, 16'd11980, 16'd26306, 16'd34975, 16'd30519, 16'd57438}; // indx = 2932
    #10;
    addra = 32'd93856;
    dina = {96'd0, 16'd54690, 16'd12889, 16'd60373, 16'd26008, 16'd23267, 16'd28910, 16'd40914, 16'd23451, 16'd13613, 16'd55956}; // indx = 2933
    #10;
    addra = 32'd93888;
    dina = {96'd0, 16'd4900, 16'd48545, 16'd1143, 16'd63297, 16'd33689, 16'd52288, 16'd54229, 16'd29037, 16'd22700, 16'd30410}; // indx = 2934
    #10;
    addra = 32'd93920;
    dina = {96'd0, 16'd31466, 16'd58678, 16'd61265, 16'd53353, 16'd65309, 16'd46573, 16'd17187, 16'd29474, 16'd61607, 16'd16815}; // indx = 2935
    #10;
    addra = 32'd93952;
    dina = {96'd0, 16'd55919, 16'd25502, 16'd17982, 16'd55806, 16'd45775, 16'd33102, 16'd32767, 16'd61238, 16'd62518, 16'd3083}; // indx = 2936
    #10;
    addra = 32'd93984;
    dina = {96'd0, 16'd23230, 16'd12758, 16'd21448, 16'd43337, 16'd17925, 16'd59407, 16'd2633, 16'd21886, 16'd22227, 16'd13652}; // indx = 2937
    #10;
    addra = 32'd94016;
    dina = {96'd0, 16'd2753, 16'd23821, 16'd28610, 16'd33076, 16'd49014, 16'd3101, 16'd59051, 16'd16454, 16'd10752, 16'd15867}; // indx = 2938
    #10;
    addra = 32'd94048;
    dina = {96'd0, 16'd50739, 16'd55428, 16'd6261, 16'd14508, 16'd29608, 16'd41734, 16'd1285, 16'd29076, 16'd44208, 16'd31940}; // indx = 2939
    #10;
    addra = 32'd94080;
    dina = {96'd0, 16'd15447, 16'd17081, 16'd9409, 16'd62898, 16'd61464, 16'd1125, 16'd58690, 16'd10633, 16'd8079, 16'd26550}; // indx = 2940
    #10;
    addra = 32'd94112;
    dina = {96'd0, 16'd31134, 16'd40594, 16'd65076, 16'd35035, 16'd24839, 16'd59933, 16'd9998, 16'd60296, 16'd64910, 16'd26950}; // indx = 2941
    #10;
    addra = 32'd94144;
    dina = {96'd0, 16'd7321, 16'd26791, 16'd61715, 16'd15652, 16'd46215, 16'd64035, 16'd22172, 16'd55007, 16'd51266, 16'd4861}; // indx = 2942
    #10;
    addra = 32'd94176;
    dina = {96'd0, 16'd21088, 16'd10509, 16'd18366, 16'd64239, 16'd4988, 16'd20474, 16'd62451, 16'd45292, 16'd42294, 16'd15843}; // indx = 2943
    #10;
    addra = 32'd94208;
    dina = {96'd0, 16'd21067, 16'd33254, 16'd26965, 16'd2238, 16'd59187, 16'd60738, 16'd3595, 16'd6859, 16'd43020, 16'd13750}; // indx = 2944
    #10;
    addra = 32'd94240;
    dina = {96'd0, 16'd26637, 16'd61067, 16'd26750, 16'd42897, 16'd44542, 16'd10527, 16'd43107, 16'd34504, 16'd46121, 16'd53039}; // indx = 2945
    #10;
    addra = 32'd94272;
    dina = {96'd0, 16'd2200, 16'd575, 16'd46658, 16'd46170, 16'd13389, 16'd65006, 16'd63637, 16'd15933, 16'd23343, 16'd13661}; // indx = 2946
    #10;
    addra = 32'd94304;
    dina = {96'd0, 16'd48649, 16'd61272, 16'd12252, 16'd57726, 16'd41960, 16'd65172, 16'd58486, 16'd51570, 16'd24658, 16'd5987}; // indx = 2947
    #10;
    addra = 32'd94336;
    dina = {96'd0, 16'd53687, 16'd29417, 16'd25179, 16'd48250, 16'd52941, 16'd27850, 16'd28473, 16'd51463, 16'd18730, 16'd63572}; // indx = 2948
    #10;
    addra = 32'd94368;
    dina = {96'd0, 16'd38695, 16'd24021, 16'd50675, 16'd37442, 16'd30092, 16'd21950, 16'd15105, 16'd8270, 16'd57549, 16'd61555}; // indx = 2949
    #10;
    addra = 32'd94400;
    dina = {96'd0, 16'd19445, 16'd30292, 16'd17766, 16'd10426, 16'd51662, 16'd32691, 16'd61179, 16'd7249, 16'd3384, 16'd34769}; // indx = 2950
    #10;
    addra = 32'd94432;
    dina = {96'd0, 16'd45055, 16'd4494, 16'd20069, 16'd62480, 16'd22152, 16'd32188, 16'd24713, 16'd62223, 16'd49832, 16'd42581}; // indx = 2951
    #10;
    addra = 32'd94464;
    dina = {96'd0, 16'd37639, 16'd57404, 16'd61402, 16'd62568, 16'd56544, 16'd18483, 16'd64884, 16'd45804, 16'd30171, 16'd5872}; // indx = 2952
    #10;
    addra = 32'd94496;
    dina = {96'd0, 16'd32181, 16'd13058, 16'd28781, 16'd27568, 16'd35227, 16'd56589, 16'd56212, 16'd7027, 16'd12238, 16'd42175}; // indx = 2953
    #10;
    addra = 32'd94528;
    dina = {96'd0, 16'd19615, 16'd42567, 16'd1526, 16'd63617, 16'd24121, 16'd19899, 16'd56968, 16'd56164, 16'd26196, 16'd57841}; // indx = 2954
    #10;
    addra = 32'd94560;
    dina = {96'd0, 16'd52006, 16'd35317, 16'd53465, 16'd30415, 16'd8633, 16'd3780, 16'd51051, 16'd64782, 16'd2723, 16'd56373}; // indx = 2955
    #10;
    addra = 32'd94592;
    dina = {96'd0, 16'd24453, 16'd39662, 16'd15188, 16'd17584, 16'd44391, 16'd49546, 16'd34076, 16'd49323, 16'd5744, 16'd32352}; // indx = 2956
    #10;
    addra = 32'd94624;
    dina = {96'd0, 16'd19289, 16'd41130, 16'd35498, 16'd43134, 16'd20484, 16'd41583, 16'd38813, 16'd40095, 16'd60141, 16'd56915}; // indx = 2957
    #10;
    addra = 32'd94656;
    dina = {96'd0, 16'd16838, 16'd57824, 16'd26109, 16'd24308, 16'd35329, 16'd27302, 16'd52325, 16'd11934, 16'd36554, 16'd25844}; // indx = 2958
    #10;
    addra = 32'd94688;
    dina = {96'd0, 16'd48641, 16'd59951, 16'd5416, 16'd7893, 16'd49170, 16'd32291, 16'd49055, 16'd49620, 16'd22496, 16'd15667}; // indx = 2959
    #10;
    addra = 32'd94720;
    dina = {96'd0, 16'd65253, 16'd16589, 16'd26651, 16'd65342, 16'd64394, 16'd600, 16'd41711, 16'd32563, 16'd31100, 16'd25396}; // indx = 2960
    #10;
    addra = 32'd94752;
    dina = {96'd0, 16'd64645, 16'd36201, 16'd5799, 16'd18676, 16'd17725, 16'd45952, 16'd49370, 16'd39169, 16'd48402, 16'd27215}; // indx = 2961
    #10;
    addra = 32'd94784;
    dina = {96'd0, 16'd61281, 16'd33696, 16'd48166, 16'd1019, 16'd26097, 16'd9581, 16'd43360, 16'd36191, 16'd21201, 16'd8241}; // indx = 2962
    #10;
    addra = 32'd94816;
    dina = {96'd0, 16'd60997, 16'd1947, 16'd9473, 16'd8297, 16'd32427, 16'd20308, 16'd65370, 16'd48949, 16'd40041, 16'd233}; // indx = 2963
    #10;
    addra = 32'd94848;
    dina = {96'd0, 16'd54365, 16'd64611, 16'd19315, 16'd38113, 16'd22954, 16'd20607, 16'd34406, 16'd5371, 16'd3816, 16'd53413}; // indx = 2964
    #10;
    addra = 32'd94880;
    dina = {96'd0, 16'd42484, 16'd11425, 16'd5177, 16'd56933, 16'd3490, 16'd62285, 16'd35255, 16'd30618, 16'd42430, 16'd43751}; // indx = 2965
    #10;
    addra = 32'd94912;
    dina = {96'd0, 16'd5072, 16'd46007, 16'd64287, 16'd38772, 16'd28322, 16'd45418, 16'd51739, 16'd26975, 16'd37638, 16'd6726}; // indx = 2966
    #10;
    addra = 32'd94944;
    dina = {96'd0, 16'd16693, 16'd23621, 16'd62537, 16'd56487, 16'd11362, 16'd5289, 16'd32485, 16'd38057, 16'd32472, 16'd47011}; // indx = 2967
    #10;
    addra = 32'd94976;
    dina = {96'd0, 16'd31068, 16'd31786, 16'd43081, 16'd21389, 16'd57283, 16'd1280, 16'd9118, 16'd2625, 16'd54291, 16'd11475}; // indx = 2968
    #10;
    addra = 32'd95008;
    dina = {96'd0, 16'd2588, 16'd19337, 16'd34745, 16'd4526, 16'd25709, 16'd8499, 16'd15816, 16'd59949, 16'd25160, 16'd12921}; // indx = 2969
    #10;
    addra = 32'd95040;
    dina = {96'd0, 16'd42567, 16'd34732, 16'd325, 16'd7214, 16'd22199, 16'd8269, 16'd9997, 16'd23211, 16'd33837, 16'd30914}; // indx = 2970
    #10;
    addra = 32'd95072;
    dina = {96'd0, 16'd143, 16'd26147, 16'd485, 16'd50534, 16'd5107, 16'd9235, 16'd26347, 16'd27671, 16'd36834, 16'd46625}; // indx = 2971
    #10;
    addra = 32'd95104;
    dina = {96'd0, 16'd20771, 16'd58158, 16'd50309, 16'd51782, 16'd30676, 16'd35494, 16'd24231, 16'd62603, 16'd57761, 16'd38809}; // indx = 2972
    #10;
    addra = 32'd95136;
    dina = {96'd0, 16'd49015, 16'd44068, 16'd63667, 16'd40354, 16'd36269, 16'd16592, 16'd1246, 16'd55403, 16'd36056, 16'd7689}; // indx = 2973
    #10;
    addra = 32'd95168;
    dina = {96'd0, 16'd49363, 16'd64395, 16'd37728, 16'd2236, 16'd21575, 16'd24843, 16'd13812, 16'd32418, 16'd16018, 16'd17904}; // indx = 2974
    #10;
    addra = 32'd95200;
    dina = {96'd0, 16'd51747, 16'd52218, 16'd64164, 16'd26503, 16'd36652, 16'd56582, 16'd8586, 16'd31039, 16'd61108, 16'd52067}; // indx = 2975
    #10;
    addra = 32'd95232;
    dina = {96'd0, 16'd5666, 16'd7169, 16'd47035, 16'd27726, 16'd20704, 16'd61143, 16'd49703, 16'd34695, 16'd4578, 16'd31249}; // indx = 2976
    #10;
    addra = 32'd95264;
    dina = {96'd0, 16'd47197, 16'd15089, 16'd31565, 16'd8688, 16'd35361, 16'd486, 16'd7074, 16'd64435, 16'd2761, 16'd11108}; // indx = 2977
    #10;
    addra = 32'd95296;
    dina = {96'd0, 16'd49726, 16'd63890, 16'd9220, 16'd29020, 16'd49598, 16'd48880, 16'd8394, 16'd20253, 16'd16019, 16'd52944}; // indx = 2978
    #10;
    addra = 32'd95328;
    dina = {96'd0, 16'd65269, 16'd42874, 16'd30609, 16'd44163, 16'd52176, 16'd47522, 16'd7599, 16'd13247, 16'd60707, 16'd32896}; // indx = 2979
    #10;
    addra = 32'd95360;
    dina = {96'd0, 16'd34864, 16'd56502, 16'd42260, 16'd18215, 16'd15069, 16'd29368, 16'd4869, 16'd64612, 16'd41228, 16'd58314}; // indx = 2980
    #10;
    addra = 32'd95392;
    dina = {96'd0, 16'd45284, 16'd36234, 16'd7467, 16'd23420, 16'd45903, 16'd43293, 16'd46812, 16'd26404, 16'd32746, 16'd46203}; // indx = 2981
    #10;
    addra = 32'd95424;
    dina = {96'd0, 16'd51657, 16'd27795, 16'd53639, 16'd41872, 16'd25168, 16'd63308, 16'd33592, 16'd43893, 16'd43607, 16'd59526}; // indx = 2982
    #10;
    addra = 32'd95456;
    dina = {96'd0, 16'd56550, 16'd9664, 16'd59848, 16'd34780, 16'd35226, 16'd2467, 16'd65416, 16'd15080, 16'd5339, 16'd35315}; // indx = 2983
    #10;
    addra = 32'd95488;
    dina = {96'd0, 16'd44993, 16'd38486, 16'd33669, 16'd38148, 16'd3206, 16'd22254, 16'd41839, 16'd35749, 16'd51487, 16'd46129}; // indx = 2984
    #10;
    addra = 32'd95520;
    dina = {96'd0, 16'd23775, 16'd20950, 16'd57968, 16'd33991, 16'd7855, 16'd42822, 16'd39867, 16'd1612, 16'd57960, 16'd40964}; // indx = 2985
    #10;
    addra = 32'd95552;
    dina = {96'd0, 16'd25236, 16'd18197, 16'd52471, 16'd26404, 16'd41901, 16'd50030, 16'd21626, 16'd42734, 16'd5389, 16'd22758}; // indx = 2986
    #10;
    addra = 32'd95584;
    dina = {96'd0, 16'd34238, 16'd31287, 16'd45684, 16'd31324, 16'd19790, 16'd43087, 16'd54092, 16'd25726, 16'd24290, 16'd22063}; // indx = 2987
    #10;
    addra = 32'd95616;
    dina = {96'd0, 16'd16955, 16'd29424, 16'd3701, 16'd63085, 16'd22926, 16'd42177, 16'd41592, 16'd21995, 16'd32313, 16'd2655}; // indx = 2988
    #10;
    addra = 32'd95648;
    dina = {96'd0, 16'd37641, 16'd7287, 16'd58781, 16'd19239, 16'd51494, 16'd44420, 16'd46450, 16'd23682, 16'd27878, 16'd17318}; // indx = 2989
    #10;
    addra = 32'd95680;
    dina = {96'd0, 16'd33606, 16'd5456, 16'd17523, 16'd34888, 16'd37539, 16'd952, 16'd6153, 16'd27179, 16'd8576, 16'd5564}; // indx = 2990
    #10;
    addra = 32'd95712;
    dina = {96'd0, 16'd39680, 16'd2968, 16'd45523, 16'd36910, 16'd12307, 16'd17691, 16'd24323, 16'd22810, 16'd13238, 16'd31018}; // indx = 2991
    #10;
    addra = 32'd95744;
    dina = {96'd0, 16'd52136, 16'd3028, 16'd27134, 16'd8079, 16'd35254, 16'd38214, 16'd19319, 16'd5066, 16'd29263, 16'd64573}; // indx = 2992
    #10;
    addra = 32'd95776;
    dina = {96'd0, 16'd10361, 16'd15281, 16'd56153, 16'd15871, 16'd32041, 16'd4129, 16'd1789, 16'd35853, 16'd5308, 16'd46168}; // indx = 2993
    #10;
    addra = 32'd95808;
    dina = {96'd0, 16'd50928, 16'd42232, 16'd11447, 16'd45532, 16'd61178, 16'd36073, 16'd52726, 16'd16989, 16'd27153, 16'd8019}; // indx = 2994
    #10;
    addra = 32'd95840;
    dina = {96'd0, 16'd7083, 16'd1373, 16'd50226, 16'd64819, 16'd63851, 16'd5646, 16'd6438, 16'd380, 16'd65390, 16'd58383}; // indx = 2995
    #10;
    addra = 32'd95872;
    dina = {96'd0, 16'd41283, 16'd15829, 16'd5260, 16'd28953, 16'd62210, 16'd17036, 16'd52246, 16'd2878, 16'd19297, 16'd61275}; // indx = 2996
    #10;
    addra = 32'd95904;
    dina = {96'd0, 16'd52875, 16'd8059, 16'd20865, 16'd46289, 16'd40749, 16'd25373, 16'd39960, 16'd34192, 16'd42257, 16'd63354}; // indx = 2997
    #10;
    addra = 32'd95936;
    dina = {96'd0, 16'd36038, 16'd39246, 16'd3250, 16'd38500, 16'd43604, 16'd45138, 16'd29502, 16'd27941, 16'd19838, 16'd20266}; // indx = 2998
    #10;
    addra = 32'd95968;
    dina = {96'd0, 16'd60319, 16'd50591, 16'd29105, 16'd47149, 16'd19863, 16'd35584, 16'd12408, 16'd30616, 16'd45307, 16'd55800}; // indx = 2999
    #10;
    addra = 32'd96000;
    dina = {96'd0, 16'd5972, 16'd17530, 16'd5356, 16'd12046, 16'd46809, 16'd13678, 16'd20366, 16'd24633, 16'd35148, 16'd41237}; // indx = 3000
    #10;
    addra = 32'd96032;
    dina = {96'd0, 16'd14282, 16'd49712, 16'd26519, 16'd59114, 16'd14132, 16'd55055, 16'd47003, 16'd61339, 16'd34460, 16'd23479}; // indx = 3001
    #10;
    addra = 32'd96064;
    dina = {96'd0, 16'd47046, 16'd40995, 16'd14978, 16'd54908, 16'd32854, 16'd47776, 16'd35166, 16'd16368, 16'd50248, 16'd11087}; // indx = 3002
    #10;
    addra = 32'd96096;
    dina = {96'd0, 16'd56578, 16'd54020, 16'd35781, 16'd13124, 16'd27396, 16'd27893, 16'd61964, 16'd63752, 16'd29640, 16'd23515}; // indx = 3003
    #10;
    addra = 32'd96128;
    dina = {96'd0, 16'd50719, 16'd11055, 16'd65375, 16'd35982, 16'd17279, 16'd10192, 16'd53255, 16'd8608, 16'd11028, 16'd50874}; // indx = 3004
    #10;
    addra = 32'd96160;
    dina = {96'd0, 16'd26961, 16'd7330, 16'd47104, 16'd36466, 16'd54500, 16'd63693, 16'd18074, 16'd35430, 16'd56469, 16'd47849}; // indx = 3005
    #10;
    addra = 32'd96192;
    dina = {96'd0, 16'd5936, 16'd15190, 16'd58809, 16'd24818, 16'd19115, 16'd34778, 16'd19919, 16'd33093, 16'd36901, 16'd19436}; // indx = 3006
    #10;
    addra = 32'd96224;
    dina = {96'd0, 16'd31607, 16'd15499, 16'd25385, 16'd50161, 16'd54661, 16'd8655, 16'd13474, 16'd38664, 16'd64648, 16'd64797}; // indx = 3007
    #10;
    addra = 32'd96256;
    dina = {96'd0, 16'd55868, 16'd16461, 16'd11221, 16'd7418, 16'd61625, 16'd14323, 16'd7614, 16'd62658, 16'd1327, 16'd32673}; // indx = 3008
    #10;
    addra = 32'd96288;
    dina = {96'd0, 16'd57502, 16'd43969, 16'd41776, 16'd41778, 16'd885, 16'd39104, 16'd41426, 16'd5672, 16'd53016, 16'd5951}; // indx = 3009
    #10;
    addra = 32'd96320;
    dina = {96'd0, 16'd9733, 16'd9809, 16'd22738, 16'd57385, 16'd52062, 16'd21029, 16'd25892, 16'd20824, 16'd13538, 16'd15219}; // indx = 3010
    #10;
    addra = 32'd96352;
    dina = {96'd0, 16'd9412, 16'd11085, 16'd14157, 16'd28517, 16'd25525, 16'd50550, 16'd44318, 16'd32863, 16'd51782, 16'd54969}; // indx = 3011
    #10;
    addra = 32'd96384;
    dina = {96'd0, 16'd61411, 16'd56322, 16'd46997, 16'd60909, 16'd5031, 16'd53643, 16'd22219, 16'd43324, 16'd38901, 16'd27615}; // indx = 3012
    #10;
    addra = 32'd96416;
    dina = {96'd0, 16'd57326, 16'd6714, 16'd3012, 16'd36884, 16'd10649, 16'd45021, 16'd57825, 16'd26725, 16'd11377, 16'd12033}; // indx = 3013
    #10;
    addra = 32'd96448;
    dina = {96'd0, 16'd19553, 16'd63387, 16'd10909, 16'd33824, 16'd40702, 16'd38167, 16'd57094, 16'd45846, 16'd12507, 16'd3085}; // indx = 3014
    #10;
    addra = 32'd96480;
    dina = {96'd0, 16'd50652, 16'd37578, 16'd19478, 16'd24877, 16'd54974, 16'd14572, 16'd9470, 16'd14770, 16'd1694, 16'd37539}; // indx = 3015
    #10;
    addra = 32'd96512;
    dina = {96'd0, 16'd51015, 16'd12060, 16'd20698, 16'd10460, 16'd21881, 16'd1044, 16'd30979, 16'd21361, 16'd19913, 16'd47220}; // indx = 3016
    #10;
    addra = 32'd96544;
    dina = {96'd0, 16'd40294, 16'd53274, 16'd7763, 16'd29045, 16'd35162, 16'd42531, 16'd20709, 16'd21525, 16'd12629, 16'd41596}; // indx = 3017
    #10;
    addra = 32'd96576;
    dina = {96'd0, 16'd11433, 16'd29096, 16'd15043, 16'd37330, 16'd25380, 16'd4673, 16'd50770, 16'd43097, 16'd21769, 16'd16726}; // indx = 3018
    #10;
    addra = 32'd96608;
    dina = {96'd0, 16'd2403, 16'd13558, 16'd8534, 16'd37738, 16'd30806, 16'd23682, 16'd16697, 16'd1954, 16'd15307, 16'd54794}; // indx = 3019
    #10;
    addra = 32'd96640;
    dina = {96'd0, 16'd432, 16'd31204, 16'd7969, 16'd52402, 16'd62727, 16'd11512, 16'd5823, 16'd51396, 16'd1794, 16'd56212}; // indx = 3020
    #10;
    addra = 32'd96672;
    dina = {96'd0, 16'd33148, 16'd16140, 16'd18153, 16'd49633, 16'd61238, 16'd46557, 16'd35171, 16'd26827, 16'd29739, 16'd65445}; // indx = 3021
    #10;
    addra = 32'd96704;
    dina = {96'd0, 16'd35772, 16'd32728, 16'd38652, 16'd12816, 16'd34195, 16'd25960, 16'd21410, 16'd9605, 16'd13487, 16'd48995}; // indx = 3022
    #10;
    addra = 32'd96736;
    dina = {96'd0, 16'd39754, 16'd6319, 16'd32905, 16'd12672, 16'd25146, 16'd42352, 16'd64406, 16'd56385, 16'd20089, 16'd39331}; // indx = 3023
    #10;
    addra = 32'd96768;
    dina = {96'd0, 16'd33968, 16'd39649, 16'd49151, 16'd31773, 16'd48690, 16'd59151, 16'd21791, 16'd22911, 16'd16474, 16'd62789}; // indx = 3024
    #10;
    addra = 32'd96800;
    dina = {96'd0, 16'd11297, 16'd65294, 16'd57002, 16'd6855, 16'd27554, 16'd31662, 16'd3508, 16'd12138, 16'd57574, 16'd15422}; // indx = 3025
    #10;
    addra = 32'd96832;
    dina = {96'd0, 16'd57789, 16'd56856, 16'd21937, 16'd16564, 16'd53822, 16'd3938, 16'd28455, 16'd3315, 16'd57181, 16'd19665}; // indx = 3026
    #10;
    addra = 32'd96864;
    dina = {96'd0, 16'd22177, 16'd11454, 16'd1644, 16'd53812, 16'd47473, 16'd39931, 16'd54940, 16'd3413, 16'd41878, 16'd32490}; // indx = 3027
    #10;
    addra = 32'd96896;
    dina = {96'd0, 16'd32090, 16'd47283, 16'd6978, 16'd38453, 16'd50899, 16'd12762, 16'd12602, 16'd39294, 16'd24391, 16'd23209}; // indx = 3028
    #10;
    addra = 32'd96928;
    dina = {96'd0, 16'd14880, 16'd47346, 16'd6550, 16'd56524, 16'd31636, 16'd38414, 16'd62867, 16'd26136, 16'd42482, 16'd45662}; // indx = 3029
    #10;
    addra = 32'd96960;
    dina = {96'd0, 16'd5414, 16'd26129, 16'd63564, 16'd38646, 16'd26834, 16'd16791, 16'd37702, 16'd56313, 16'd7246, 16'd45946}; // indx = 3030
    #10;
    addra = 32'd96992;
    dina = {96'd0, 16'd51, 16'd28850, 16'd56989, 16'd56226, 16'd65084, 16'd13938, 16'd63726, 16'd16296, 16'd52380, 16'd40367}; // indx = 3031
    #10;
    addra = 32'd97024;
    dina = {96'd0, 16'd14002, 16'd21201, 16'd5420, 16'd64895, 16'd3177, 16'd43894, 16'd62336, 16'd39502, 16'd22766, 16'd44387}; // indx = 3032
    #10;
    addra = 32'd97056;
    dina = {96'd0, 16'd33696, 16'd21589, 16'd41109, 16'd3891, 16'd28916, 16'd8812, 16'd11733, 16'd47125, 16'd21759, 16'd65082}; // indx = 3033
    #10;
    addra = 32'd97088;
    dina = {96'd0, 16'd58280, 16'd13548, 16'd33330, 16'd8594, 16'd8387, 16'd22989, 16'd50948, 16'd56106, 16'd61185, 16'd41905}; // indx = 3034
    #10;
    addra = 32'd97120;
    dina = {96'd0, 16'd5311, 16'd58813, 16'd45840, 16'd20429, 16'd10488, 16'd374, 16'd33723, 16'd59177, 16'd58573, 16'd346}; // indx = 3035
    #10;
    addra = 32'd97152;
    dina = {96'd0, 16'd50468, 16'd45211, 16'd41969, 16'd62342, 16'd45898, 16'd11922, 16'd18366, 16'd2307, 16'd41357, 16'd57151}; // indx = 3036
    #10;
    addra = 32'd97184;
    dina = {96'd0, 16'd63123, 16'd39062, 16'd53790, 16'd18485, 16'd35467, 16'd50567, 16'd58194, 16'd23904, 16'd23325, 16'd19242}; // indx = 3037
    #10;
    addra = 32'd97216;
    dina = {96'd0, 16'd5273, 16'd62224, 16'd21478, 16'd63764, 16'd12071, 16'd57463, 16'd25412, 16'd37805, 16'd19596, 16'd19556}; // indx = 3038
    #10;
    addra = 32'd97248;
    dina = {96'd0, 16'd1635, 16'd44074, 16'd16701, 16'd56919, 16'd40479, 16'd44635, 16'd3676, 16'd24864, 16'd32357, 16'd2170}; // indx = 3039
    #10;
    addra = 32'd97280;
    dina = {96'd0, 16'd30581, 16'd35925, 16'd46794, 16'd48901, 16'd14594, 16'd55482, 16'd41317, 16'd42129, 16'd8145, 16'd29408}; // indx = 3040
    #10;
    addra = 32'd97312;
    dina = {96'd0, 16'd7883, 16'd63388, 16'd21728, 16'd56811, 16'd26598, 16'd6819, 16'd11679, 16'd11694, 16'd47130, 16'd9465}; // indx = 3041
    #10;
    addra = 32'd97344;
    dina = {96'd0, 16'd46805, 16'd19643, 16'd9064, 16'd26242, 16'd46828, 16'd19073, 16'd39026, 16'd28916, 16'd20520, 16'd24954}; // indx = 3042
    #10;
    addra = 32'd97376;
    dina = {96'd0, 16'd47419, 16'd62940, 16'd41325, 16'd6779, 16'd41607, 16'd15058, 16'd18816, 16'd48367, 16'd45858, 16'd29851}; // indx = 3043
    #10;
    addra = 32'd97408;
    dina = {96'd0, 16'd57365, 16'd56874, 16'd20184, 16'd31618, 16'd23519, 16'd64979, 16'd37832, 16'd7212, 16'd43734, 16'd26465}; // indx = 3044
    #10;
    addra = 32'd97440;
    dina = {96'd0, 16'd38966, 16'd16613, 16'd16584, 16'd22056, 16'd13960, 16'd56666, 16'd31760, 16'd17923, 16'd55585, 16'd33617}; // indx = 3045
    #10;
    addra = 32'd97472;
    dina = {96'd0, 16'd53908, 16'd2662, 16'd47783, 16'd12841, 16'd17821, 16'd11467, 16'd60819, 16'd34606, 16'd13365, 16'd59829}; // indx = 3046
    #10;
    addra = 32'd97504;
    dina = {96'd0, 16'd53851, 16'd1345, 16'd39648, 16'd36450, 16'd35726, 16'd2373, 16'd21557, 16'd26162, 16'd35848, 16'd51691}; // indx = 3047
    #10;
    addra = 32'd97536;
    dina = {96'd0, 16'd40448, 16'd32534, 16'd2210, 16'd16950, 16'd8611, 16'd35515, 16'd35652, 16'd65113, 16'd32648, 16'd42361}; // indx = 3048
    #10;
    addra = 32'd97568;
    dina = {96'd0, 16'd12517, 16'd14402, 16'd22260, 16'd43137, 16'd36900, 16'd60559, 16'd65304, 16'd29526, 16'd16074, 16'd48458}; // indx = 3049
    #10;
    addra = 32'd97600;
    dina = {96'd0, 16'd12591, 16'd24243, 16'd32961, 16'd7897, 16'd64199, 16'd2367, 16'd1052, 16'd10262, 16'd27257, 16'd11194}; // indx = 3050
    #10;
    addra = 32'd97632;
    dina = {96'd0, 16'd49177, 16'd50562, 16'd31905, 16'd31846, 16'd54919, 16'd1002, 16'd44369, 16'd30813, 16'd64722, 16'd59409}; // indx = 3051
    #10;
    addra = 32'd97664;
    dina = {96'd0, 16'd11167, 16'd24206, 16'd49180, 16'd39327, 16'd27981, 16'd24182, 16'd46146, 16'd26148, 16'd6836, 16'd31347}; // indx = 3052
    #10;
    addra = 32'd97696;
    dina = {96'd0, 16'd14545, 16'd60431, 16'd26076, 16'd32455, 16'd2558, 16'd27880, 16'd1720, 16'd40746, 16'd8750, 16'd10796}; // indx = 3053
    #10;
    addra = 32'd97728;
    dina = {96'd0, 16'd49370, 16'd58655, 16'd25885, 16'd43821, 16'd9542, 16'd47732, 16'd52776, 16'd17746, 16'd35337, 16'd29837}; // indx = 3054
    #10;
    addra = 32'd97760;
    dina = {96'd0, 16'd39879, 16'd46787, 16'd57424, 16'd14510, 16'd53707, 16'd44655, 16'd36055, 16'd22152, 16'd54018, 16'd17961}; // indx = 3055
    #10;
    addra = 32'd97792;
    dina = {96'd0, 16'd5858, 16'd43086, 16'd29422, 16'd39786, 16'd26604, 16'd44952, 16'd59851, 16'd14945, 16'd58536, 16'd26689}; // indx = 3056
    #10;
    addra = 32'd97824;
    dina = {96'd0, 16'd45333, 16'd34431, 16'd12847, 16'd42597, 16'd31029, 16'd39933, 16'd38043, 16'd9543, 16'd8468, 16'd33711}; // indx = 3057
    #10;
    addra = 32'd97856;
    dina = {96'd0, 16'd19616, 16'd29863, 16'd36656, 16'd18485, 16'd54307, 16'd41565, 16'd30995, 16'd4339, 16'd51111, 16'd36115}; // indx = 3058
    #10;
    addra = 32'd97888;
    dina = {96'd0, 16'd8280, 16'd19497, 16'd48780, 16'd33546, 16'd27118, 16'd40399, 16'd15630, 16'd14809, 16'd25512, 16'd21823}; // indx = 3059
    #10;
    addra = 32'd97920;
    dina = {96'd0, 16'd20019, 16'd35333, 16'd31873, 16'd18994, 16'd675, 16'd43627, 16'd55339, 16'd27625, 16'd7917, 16'd52603}; // indx = 3060
    #10;
    addra = 32'd97952;
    dina = {96'd0, 16'd23233, 16'd32575, 16'd60917, 16'd13182, 16'd50450, 16'd12938, 16'd65240, 16'd50303, 16'd20310, 16'd37405}; // indx = 3061
    #10;
    addra = 32'd97984;
    dina = {96'd0, 16'd11805, 16'd43870, 16'd5051, 16'd50865, 16'd21526, 16'd41580, 16'd47871, 16'd28517, 16'd24782, 16'd18700}; // indx = 3062
    #10;
    addra = 32'd98016;
    dina = {96'd0, 16'd29542, 16'd44075, 16'd38046, 16'd35334, 16'd36576, 16'd33974, 16'd59361, 16'd59596, 16'd39849, 16'd53323}; // indx = 3063
    #10;
    addra = 32'd98048;
    dina = {96'd0, 16'd18828, 16'd43297, 16'd10175, 16'd10752, 16'd30093, 16'd42115, 16'd41598, 16'd26046, 16'd15962, 16'd11304}; // indx = 3064
    #10;
    addra = 32'd98080;
    dina = {96'd0, 16'd36985, 16'd26804, 16'd43688, 16'd13753, 16'd5589, 16'd11048, 16'd14270, 16'd11502, 16'd52845, 16'd56008}; // indx = 3065
    #10;
    addra = 32'd98112;
    dina = {96'd0, 16'd13263, 16'd33430, 16'd33713, 16'd22877, 16'd31843, 16'd61742, 16'd62672, 16'd32222, 16'd53603, 16'd56371}; // indx = 3066
    #10;
    addra = 32'd98144;
    dina = {96'd0, 16'd21125, 16'd19003, 16'd23364, 16'd17801, 16'd6180, 16'd36351, 16'd51765, 16'd42612, 16'd59625, 16'd55179}; // indx = 3067
    #10;
    addra = 32'd98176;
    dina = {96'd0, 16'd60234, 16'd20221, 16'd5134, 16'd46809, 16'd27475, 16'd6087, 16'd62204, 16'd9483, 16'd10272, 16'd19719}; // indx = 3068
    #10;
    addra = 32'd98208;
    dina = {96'd0, 16'd6408, 16'd35683, 16'd27231, 16'd18337, 16'd57075, 16'd31055, 16'd16439, 16'd26372, 16'd10116, 16'd53119}; // indx = 3069
    #10;
    addra = 32'd98240;
    dina = {96'd0, 16'd4663, 16'd47561, 16'd24392, 16'd8915, 16'd63840, 16'd55613, 16'd15884, 16'd64372, 16'd57852, 16'd19722}; // indx = 3070
    #10;
    addra = 32'd98272;
    dina = {96'd0, 16'd41704, 16'd34366, 16'd54167, 16'd42370, 16'd19721, 16'd53709, 16'd28740, 16'd43458, 16'd14535, 16'd15243}; // indx = 3071
    #10;
    addra = 32'd98304;
    dina = {96'd0, 16'd6385, 16'd38228, 16'd30091, 16'd60524, 16'd54258, 16'd53210, 16'd59110, 16'd35462, 16'd18319, 16'd20012}; // indx = 3072
    #10;
    addra = 32'd98336;
    dina = {96'd0, 16'd42600, 16'd29445, 16'd16711, 16'd39788, 16'd32980, 16'd5939, 16'd45850, 16'd60735, 16'd59298, 16'd11980}; // indx = 3073
    #10;
    addra = 32'd98368;
    dina = {96'd0, 16'd50656, 16'd19622, 16'd13298, 16'd51145, 16'd21353, 16'd20469, 16'd34075, 16'd23131, 16'd7657, 16'd57130}; // indx = 3074
    #10;
    addra = 32'd98400;
    dina = {96'd0, 16'd32230, 16'd20857, 16'd46580, 16'd57701, 16'd63181, 16'd44325, 16'd61794, 16'd50911, 16'd19323, 16'd40498}; // indx = 3075
    #10;
    addra = 32'd98432;
    dina = {96'd0, 16'd36304, 16'd47060, 16'd60328, 16'd31393, 16'd45917, 16'd52150, 16'd11028, 16'd29854, 16'd28709, 16'd32020}; // indx = 3076
    #10;
    addra = 32'd98464;
    dina = {96'd0, 16'd51191, 16'd18544, 16'd11982, 16'd11292, 16'd57398, 16'd16788, 16'd19221, 16'd69, 16'd37885, 16'd35325}; // indx = 3077
    #10;
    addra = 32'd98496;
    dina = {96'd0, 16'd20978, 16'd65170, 16'd39137, 16'd9778, 16'd62803, 16'd59056, 16'd61794, 16'd43560, 16'd18622, 16'd18131}; // indx = 3078
    #10;
    addra = 32'd98528;
    dina = {96'd0, 16'd32444, 16'd27245, 16'd60148, 16'd19794, 16'd44955, 16'd31036, 16'd14029, 16'd51018, 16'd65252, 16'd7317}; // indx = 3079
    #10;
    addra = 32'd98560;
    dina = {96'd0, 16'd5203, 16'd28122, 16'd64836, 16'd54555, 16'd17303, 16'd29722, 16'd34470, 16'd3010, 16'd51882, 16'd63112}; // indx = 3080
    #10;
    addra = 32'd98592;
    dina = {96'd0, 16'd2194, 16'd41468, 16'd58756, 16'd54006, 16'd13478, 16'd30900, 16'd19681, 16'd47948, 16'd27656, 16'd40791}; // indx = 3081
    #10;
    addra = 32'd98624;
    dina = {96'd0, 16'd59925, 16'd53988, 16'd4810, 16'd34255, 16'd11047, 16'd51180, 16'd18448, 16'd6824, 16'd63772, 16'd51491}; // indx = 3082
    #10;
    addra = 32'd98656;
    dina = {96'd0, 16'd22931, 16'd12155, 16'd25224, 16'd30404, 16'd4532, 16'd27124, 16'd17361, 16'd65484, 16'd48227, 16'd36727}; // indx = 3083
    #10;
    addra = 32'd98688;
    dina = {96'd0, 16'd13919, 16'd17920, 16'd19071, 16'd19323, 16'd62131, 16'd55566, 16'd49603, 16'd56925, 16'd8453, 16'd20675}; // indx = 3084
    #10;
    addra = 32'd98720;
    dina = {96'd0, 16'd26170, 16'd39573, 16'd61746, 16'd30991, 16'd60096, 16'd826, 16'd35775, 16'd30241, 16'd18578, 16'd10535}; // indx = 3085
    #10;
    addra = 32'd98752;
    dina = {96'd0, 16'd25434, 16'd23124, 16'd15192, 16'd6154, 16'd63688, 16'd21256, 16'd23580, 16'd48829, 16'd1610, 16'd46064}; // indx = 3086
    #10;
    addra = 32'd98784;
    dina = {96'd0, 16'd45979, 16'd55051, 16'd57976, 16'd59876, 16'd50498, 16'd43565, 16'd40533, 16'd53612, 16'd63118, 16'd18336}; // indx = 3087
    #10;
    addra = 32'd98816;
    dina = {96'd0, 16'd24836, 16'd43543, 16'd29555, 16'd1649, 16'd41603, 16'd16299, 16'd59511, 16'd64309, 16'd2524, 16'd1642}; // indx = 3088
    #10;
    addra = 32'd98848;
    dina = {96'd0, 16'd49001, 16'd61718, 16'd22582, 16'd47805, 16'd43065, 16'd37538, 16'd486, 16'd28213, 16'd51235, 16'd41068}; // indx = 3089
    #10;
    addra = 32'd98880;
    dina = {96'd0, 16'd54935, 16'd47423, 16'd2149, 16'd5223, 16'd40952, 16'd9344, 16'd30091, 16'd39286, 16'd56199, 16'd23968}; // indx = 3090
    #10;
    addra = 32'd98912;
    dina = {96'd0, 16'd18314, 16'd56428, 16'd4439, 16'd54378, 16'd63229, 16'd10318, 16'd63728, 16'd55222, 16'd22982, 16'd34183}; // indx = 3091
    #10;
    addra = 32'd98944;
    dina = {96'd0, 16'd47705, 16'd942, 16'd8498, 16'd21347, 16'd37692, 16'd42940, 16'd31605, 16'd56844, 16'd54049, 16'd10979}; // indx = 3092
    #10;
    addra = 32'd98976;
    dina = {96'd0, 16'd61199, 16'd4017, 16'd3488, 16'd57620, 16'd11623, 16'd20541, 16'd42173, 16'd18822, 16'd56302, 16'd11921}; // indx = 3093
    #10;
    addra = 32'd99008;
    dina = {96'd0, 16'd64511, 16'd29392, 16'd52571, 16'd28568, 16'd60486, 16'd20874, 16'd56061, 16'd43789, 16'd37030, 16'd32740}; // indx = 3094
    #10;
    addra = 32'd99040;
    dina = {96'd0, 16'd43159, 16'd64827, 16'd59405, 16'd23798, 16'd45730, 16'd48685, 16'd18054, 16'd35417, 16'd62618, 16'd34287}; // indx = 3095
    #10;
    addra = 32'd99072;
    dina = {96'd0, 16'd5018, 16'd39141, 16'd5704, 16'd44281, 16'd2189, 16'd9411, 16'd63937, 16'd36983, 16'd62609, 16'd44573}; // indx = 3096
    #10;
    addra = 32'd99104;
    dina = {96'd0, 16'd53552, 16'd31239, 16'd49075, 16'd63776, 16'd41582, 16'd47584, 16'd12100, 16'd43630, 16'd3900, 16'd430}; // indx = 3097
    #10;
    addra = 32'd99136;
    dina = {96'd0, 16'd2133, 16'd51941, 16'd53466, 16'd29454, 16'd54154, 16'd44765, 16'd57358, 16'd64572, 16'd62479, 16'd30125}; // indx = 3098
    #10;
    addra = 32'd99168;
    dina = {96'd0, 16'd64685, 16'd50720, 16'd41679, 16'd38079, 16'd27783, 16'd21964, 16'd3347, 16'd22419, 16'd57379, 16'd25175}; // indx = 3099
    #10;
    addra = 32'd99200;
    dina = {96'd0, 16'd38708, 16'd39641, 16'd45453, 16'd56523, 16'd44269, 16'd45529, 16'd24784, 16'd60031, 16'd54876, 16'd34015}; // indx = 3100
    #10;
    addra = 32'd99232;
    dina = {96'd0, 16'd48150, 16'd33850, 16'd50621, 16'd13160, 16'd21604, 16'd10418, 16'd30732, 16'd21648, 16'd1053, 16'd47760}; // indx = 3101
    #10;
    addra = 32'd99264;
    dina = {96'd0, 16'd63687, 16'd38951, 16'd40301, 16'd18919, 16'd58826, 16'd29101, 16'd64396, 16'd40062, 16'd64360, 16'd16760}; // indx = 3102
    #10;
    addra = 32'd99296;
    dina = {96'd0, 16'd64537, 16'd33549, 16'd64927, 16'd19984, 16'd6501, 16'd31089, 16'd43549, 16'd22863, 16'd64953, 16'd23218}; // indx = 3103
    #10;
    addra = 32'd99328;
    dina = {96'd0, 16'd5026, 16'd18296, 16'd13485, 16'd20787, 16'd17969, 16'd58063, 16'd48658, 16'd4911, 16'd5747, 16'd9075}; // indx = 3104
    #10;
    addra = 32'd99360;
    dina = {96'd0, 16'd21310, 16'd47289, 16'd50760, 16'd57982, 16'd29627, 16'd52443, 16'd57722, 16'd14600, 16'd57957, 16'd51140}; // indx = 3105
    #10;
    addra = 32'd99392;
    dina = {96'd0, 16'd62197, 16'd47386, 16'd15910, 16'd38201, 16'd17012, 16'd52627, 16'd38209, 16'd17216, 16'd35227, 16'd24097}; // indx = 3106
    #10;
    addra = 32'd99424;
    dina = {96'd0, 16'd12114, 16'd24885, 16'd20468, 16'd40512, 16'd42872, 16'd11773, 16'd56974, 16'd10851, 16'd2179, 16'd20841}; // indx = 3107
    #10;
    addra = 32'd99456;
    dina = {96'd0, 16'd45802, 16'd54233, 16'd16164, 16'd63570, 16'd32899, 16'd58484, 16'd39852, 16'd48085, 16'd9245, 16'd20797}; // indx = 3108
    #10;
    addra = 32'd99488;
    dina = {96'd0, 16'd42532, 16'd16782, 16'd42682, 16'd15200, 16'd3901, 16'd2702, 16'd26078, 16'd36554, 16'd3167, 16'd42748}; // indx = 3109
    #10;
    addra = 32'd99520;
    dina = {96'd0, 16'd38794, 16'd10113, 16'd31510, 16'd21029, 16'd62488, 16'd5174, 16'd3633, 16'd65016, 16'd53282, 16'd23353}; // indx = 3110
    #10;
    addra = 32'd99552;
    dina = {96'd0, 16'd60342, 16'd40093, 16'd45459, 16'd63362, 16'd54254, 16'd29044, 16'd30758, 16'd36708, 16'd4956, 16'd34171}; // indx = 3111
    #10;
    addra = 32'd99584;
    dina = {96'd0, 16'd8293, 16'd41967, 16'd55401, 16'd21149, 16'd19208, 16'd6826, 16'd19482, 16'd21230, 16'd54205, 16'd19280}; // indx = 3112
    #10;
    addra = 32'd99616;
    dina = {96'd0, 16'd53915, 16'd18433, 16'd43354, 16'd61033, 16'd65503, 16'd8042, 16'd53898, 16'd64454, 16'd56002, 16'd41126}; // indx = 3113
    #10;
    addra = 32'd99648;
    dina = {96'd0, 16'd53992, 16'd36183, 16'd50578, 16'd7052, 16'd26411, 16'd54851, 16'd9274, 16'd47583, 16'd51455, 16'd32170}; // indx = 3114
    #10;
    addra = 32'd99680;
    dina = {96'd0, 16'd24179, 16'd23024, 16'd54660, 16'd2585, 16'd10521, 16'd52507, 16'd9068, 16'd50743, 16'd64254, 16'd35536}; // indx = 3115
    #10;
    addra = 32'd99712;
    dina = {96'd0, 16'd59536, 16'd53799, 16'd24228, 16'd40682, 16'd27571, 16'd52817, 16'd36754, 16'd23096, 16'd22974, 16'd38002}; // indx = 3116
    #10;
    addra = 32'd99744;
    dina = {96'd0, 16'd47610, 16'd566, 16'd58714, 16'd51333, 16'd44386, 16'd22047, 16'd44666, 16'd8917, 16'd28511, 16'd15877}; // indx = 3117
    #10;
    addra = 32'd99776;
    dina = {96'd0, 16'd6842, 16'd9182, 16'd32770, 16'd20450, 16'd49810, 16'd48117, 16'd60241, 16'd26747, 16'd25755, 16'd52067}; // indx = 3118
    #10;
    addra = 32'd99808;
    dina = {96'd0, 16'd12229, 16'd21785, 16'd19506, 16'd63569, 16'd44270, 16'd19914, 16'd12314, 16'd51292, 16'd13219, 16'd49712}; // indx = 3119
    #10;
    addra = 32'd99840;
    dina = {96'd0, 16'd34347, 16'd19073, 16'd64105, 16'd2000, 16'd46887, 16'd38788, 16'd1922, 16'd43057, 16'd12927, 16'd49960}; // indx = 3120
    #10;
    addra = 32'd99872;
    dina = {96'd0, 16'd2710, 16'd53722, 16'd25108, 16'd59744, 16'd60353, 16'd39364, 16'd3926, 16'd36551, 16'd1264, 16'd499}; // indx = 3121
    #10;
    addra = 32'd99904;
    dina = {96'd0, 16'd46777, 16'd12581, 16'd31287, 16'd51350, 16'd14863, 16'd11282, 16'd32070, 16'd43123, 16'd49748, 16'd15518}; // indx = 3122
    #10;
    addra = 32'd99936;
    dina = {96'd0, 16'd44358, 16'd56647, 16'd48717, 16'd52831, 16'd9009, 16'd28930, 16'd65376, 16'd31313, 16'd26335, 16'd18850}; // indx = 3123
    #10;
    addra = 32'd99968;
    dina = {96'd0, 16'd3713, 16'd11014, 16'd12250, 16'd36228, 16'd42138, 16'd5938, 16'd63849, 16'd60103, 16'd38840, 16'd38478}; // indx = 3124
    #10;
    addra = 32'd100000;
    dina = {96'd0, 16'd35304, 16'd62518, 16'd9695, 16'd13692, 16'd21472, 16'd26527, 16'd8487, 16'd47107, 16'd39527, 16'd56095}; // indx = 3125
    #10;
    addra = 32'd100032;
    dina = {96'd0, 16'd34597, 16'd44094, 16'd47391, 16'd17020, 16'd33040, 16'd10560, 16'd54517, 16'd23100, 16'd42296, 16'd1729}; // indx = 3126
    #10;
    addra = 32'd100064;
    dina = {96'd0, 16'd45750, 16'd22989, 16'd19426, 16'd12240, 16'd6716, 16'd18979, 16'd23810, 16'd57056, 16'd23536, 16'd62396}; // indx = 3127
    #10;
    addra = 32'd100096;
    dina = {96'd0, 16'd3278, 16'd33251, 16'd6730, 16'd30196, 16'd30582, 16'd27042, 16'd55995, 16'd45945, 16'd63415, 16'd43630}; // indx = 3128
    #10;
    addra = 32'd100128;
    dina = {96'd0, 16'd46689, 16'd47751, 16'd46538, 16'd58657, 16'd7019, 16'd12548, 16'd65416, 16'd64012, 16'd15817, 16'd8758}; // indx = 3129
    #10;
    addra = 32'd100160;
    dina = {96'd0, 16'd29073, 16'd11516, 16'd53826, 16'd8470, 16'd63544, 16'd64733, 16'd24487, 16'd28573, 16'd43150, 16'd25613}; // indx = 3130
    #10;
    addra = 32'd100192;
    dina = {96'd0, 16'd13533, 16'd54567, 16'd3287, 16'd3889, 16'd57629, 16'd8237, 16'd57563, 16'd63177, 16'd40711, 16'd26411}; // indx = 3131
    #10;
    addra = 32'd100224;
    dina = {96'd0, 16'd61741, 16'd32003, 16'd18799, 16'd29371, 16'd28848, 16'd44066, 16'd33780, 16'd25966, 16'd1207, 16'd46954}; // indx = 3132
    #10;
    addra = 32'd100256;
    dina = {96'd0, 16'd59950, 16'd43771, 16'd22192, 16'd42818, 16'd32448, 16'd16234, 16'd50906, 16'd33686, 16'd65107, 16'd37587}; // indx = 3133
    #10;
    addra = 32'd100288;
    dina = {96'd0, 16'd60185, 16'd42133, 16'd9848, 16'd58075, 16'd51750, 16'd15096, 16'd47706, 16'd43129, 16'd39625, 16'd22605}; // indx = 3134
    #10;
    addra = 32'd100320;
    dina = {96'd0, 16'd27318, 16'd9925, 16'd1099, 16'd6672, 16'd9384, 16'd39338, 16'd520, 16'd22039, 16'd37752, 16'd3469}; // indx = 3135
    #10;
    addra = 32'd100352;
    dina = {96'd0, 16'd25699, 16'd24847, 16'd9121, 16'd26881, 16'd39160, 16'd53784, 16'd61404, 16'd415, 16'd48626, 16'd10722}; // indx = 3136
    #10;
    addra = 32'd100384;
    dina = {96'd0, 16'd28478, 16'd61996, 16'd43001, 16'd25961, 16'd46092, 16'd20289, 16'd18992, 16'd46472, 16'd61828, 16'd49837}; // indx = 3137
    #10;
    addra = 32'd100416;
    dina = {96'd0, 16'd61812, 16'd58541, 16'd60379, 16'd3257, 16'd48051, 16'd3591, 16'd65208, 16'd32578, 16'd62351, 16'd27584}; // indx = 3138
    #10;
    addra = 32'd100448;
    dina = {96'd0, 16'd47595, 16'd61629, 16'd39333, 16'd60072, 16'd2975, 16'd25865, 16'd52135, 16'd43650, 16'd1958, 16'd44291}; // indx = 3139
    #10;
    addra = 32'd100480;
    dina = {96'd0, 16'd42957, 16'd34919, 16'd65466, 16'd10179, 16'd56556, 16'd10942, 16'd23531, 16'd21977, 16'd26684, 16'd49914}; // indx = 3140
    #10;
    addra = 32'd100512;
    dina = {96'd0, 16'd62007, 16'd17130, 16'd42335, 16'd26918, 16'd47949, 16'd18866, 16'd3692, 16'd58182, 16'd18133, 16'd51410}; // indx = 3141
    #10;
    addra = 32'd100544;
    dina = {96'd0, 16'd62796, 16'd19535, 16'd41432, 16'd57571, 16'd13110, 16'd63301, 16'd62778, 16'd48192, 16'd57275, 16'd16386}; // indx = 3142
    #10;
    addra = 32'd100576;
    dina = {96'd0, 16'd59466, 16'd48750, 16'd45813, 16'd15579, 16'd9970, 16'd24574, 16'd50269, 16'd13213, 16'd49156, 16'd55997}; // indx = 3143
    #10;
    addra = 32'd100608;
    dina = {96'd0, 16'd25752, 16'd24109, 16'd35328, 16'd40972, 16'd56044, 16'd59439, 16'd9052, 16'd44983, 16'd13124, 16'd48137}; // indx = 3144
    #10;
    addra = 32'd100640;
    dina = {96'd0, 16'd33309, 16'd60116, 16'd41525, 16'd26972, 16'd6403, 16'd28492, 16'd41920, 16'd8970, 16'd64590, 16'd30286}; // indx = 3145
    #10;
    addra = 32'd100672;
    dina = {96'd0, 16'd60893, 16'd34138, 16'd38625, 16'd59973, 16'd40834, 16'd5872, 16'd20489, 16'd37073, 16'd43930, 16'd57093}; // indx = 3146
    #10;
    addra = 32'd100704;
    dina = {96'd0, 16'd31402, 16'd22308, 16'd63957, 16'd21509, 16'd34491, 16'd18213, 16'd59600, 16'd5304, 16'd33976, 16'd23410}; // indx = 3147
    #10;
    addra = 32'd100736;
    dina = {96'd0, 16'd17867, 16'd8714, 16'd10223, 16'd4254, 16'd24038, 16'd40359, 16'd50679, 16'd1402, 16'd1871, 16'd39134}; // indx = 3148
    #10;
    addra = 32'd100768;
    dina = {96'd0, 16'd30466, 16'd17394, 16'd47871, 16'd44195, 16'd65379, 16'd14774, 16'd12244, 16'd63265, 16'd54738, 16'd37006}; // indx = 3149
    #10;
    addra = 32'd100800;
    dina = {96'd0, 16'd19007, 16'd55864, 16'd12619, 16'd31058, 16'd4757, 16'd51261, 16'd49986, 16'd17671, 16'd2648, 16'd16760}; // indx = 3150
    #10;
    addra = 32'd100832;
    dina = {96'd0, 16'd11261, 16'd37294, 16'd1936, 16'd25201, 16'd45470, 16'd41811, 16'd2249, 16'd60177, 16'd20391, 16'd8143}; // indx = 3151
    #10;
    addra = 32'd100864;
    dina = {96'd0, 16'd40126, 16'd9456, 16'd44999, 16'd40686, 16'd35070, 16'd46991, 16'd7858, 16'd48555, 16'd27883, 16'd64459}; // indx = 3152
    #10;
    addra = 32'd100896;
    dina = {96'd0, 16'd44788, 16'd56243, 16'd25809, 16'd61869, 16'd43958, 16'd53466, 16'd43586, 16'd58202, 16'd14391, 16'd53379}; // indx = 3153
    #10;
    addra = 32'd100928;
    dina = {96'd0, 16'd40244, 16'd33234, 16'd30283, 16'd58115, 16'd46339, 16'd43310, 16'd8671, 16'd35933, 16'd25005, 16'd8159}; // indx = 3154
    #10;
    addra = 32'd100960;
    dina = {96'd0, 16'd49669, 16'd35770, 16'd26587, 16'd48132, 16'd7210, 16'd12922, 16'd61928, 16'd58560, 16'd64758, 16'd30341}; // indx = 3155
    #10;
    addra = 32'd100992;
    dina = {96'd0, 16'd10384, 16'd10989, 16'd19943, 16'd38438, 16'd5690, 16'd48529, 16'd31725, 16'd34746, 16'd63389, 16'd1352}; // indx = 3156
    #10;
    addra = 32'd101024;
    dina = {96'd0, 16'd38018, 16'd62200, 16'd42002, 16'd3035, 16'd20603, 16'd29791, 16'd39471, 16'd43115, 16'd61250, 16'd51560}; // indx = 3157
    #10;
    addra = 32'd101056;
    dina = {96'd0, 16'd30178, 16'd12101, 16'd9260, 16'd52198, 16'd52725, 16'd49356, 16'd47273, 16'd8136, 16'd45169, 16'd27917}; // indx = 3158
    #10;
    addra = 32'd101088;
    dina = {96'd0, 16'd36506, 16'd36643, 16'd51779, 16'd32764, 16'd45219, 16'd25226, 16'd9734, 16'd11435, 16'd59059, 16'd35743}; // indx = 3159
    #10;
    addra = 32'd101120;
    dina = {96'd0, 16'd3119, 16'd17813, 16'd10003, 16'd55299, 16'd5557, 16'd1235, 16'd55621, 16'd28489, 16'd37724, 16'd27947}; // indx = 3160
    #10;
    addra = 32'd101152;
    dina = {96'd0, 16'd60435, 16'd64967, 16'd2385, 16'd12228, 16'd43288, 16'd14083, 16'd38676, 16'd25383, 16'd34039, 16'd12925}; // indx = 3161
    #10;
    addra = 32'd101184;
    dina = {96'd0, 16'd29509, 16'd477, 16'd23443, 16'd16702, 16'd12366, 16'd6771, 16'd58634, 16'd10324, 16'd1823, 16'd60837}; // indx = 3162
    #10;
    addra = 32'd101216;
    dina = {96'd0, 16'd24239, 16'd59616, 16'd13697, 16'd7264, 16'd40943, 16'd58296, 16'd18744, 16'd19423, 16'd22457, 16'd38341}; // indx = 3163
    #10;
    addra = 32'd101248;
    dina = {96'd0, 16'd56908, 16'd36586, 16'd35046, 16'd58945, 16'd2212, 16'd4770, 16'd25294, 16'd56882, 16'd47477, 16'd51793}; // indx = 3164
    #10;
    addra = 32'd101280;
    dina = {96'd0, 16'd50534, 16'd7039, 16'd62051, 16'd50327, 16'd10220, 16'd50357, 16'd49773, 16'd45261, 16'd14659, 16'd23498}; // indx = 3165
    #10;
    addra = 32'd101312;
    dina = {96'd0, 16'd59591, 16'd53708, 16'd20233, 16'd7143, 16'd55790, 16'd2498, 16'd36920, 16'd33458, 16'd29847, 16'd50382}; // indx = 3166
    #10;
    addra = 32'd101344;
    dina = {96'd0, 16'd63915, 16'd51631, 16'd22838, 16'd1065, 16'd39907, 16'd17355, 16'd57511, 16'd24943, 16'd39669, 16'd11308}; // indx = 3167
    #10;
    addra = 32'd101376;
    dina = {96'd0, 16'd39563, 16'd45199, 16'd2294, 16'd45368, 16'd25084, 16'd38480, 16'd61753, 16'd40672, 16'd36888, 16'd63411}; // indx = 3168
    #10;
    addra = 32'd101408;
    dina = {96'd0, 16'd16175, 16'd40940, 16'd1806, 16'd21298, 16'd16427, 16'd39371, 16'd50481, 16'd6674, 16'd38695, 16'd63982}; // indx = 3169
    #10;
    addra = 32'd101440;
    dina = {96'd0, 16'd24084, 16'd31336, 16'd57982, 16'd14196, 16'd9479, 16'd20599, 16'd58660, 16'd43498, 16'd47892, 16'd1491}; // indx = 3170
    #10;
    addra = 32'd101472;
    dina = {96'd0, 16'd11906, 16'd1017, 16'd34600, 16'd32866, 16'd38566, 16'd34567, 16'd23676, 16'd47892, 16'd10557, 16'd15283}; // indx = 3171
    #10;
    addra = 32'd101504;
    dina = {96'd0, 16'd27647, 16'd28870, 16'd32922, 16'd16396, 16'd16203, 16'd28866, 16'd34774, 16'd57707, 16'd4083, 16'd42087}; // indx = 3172
    #10;
    addra = 32'd101536;
    dina = {96'd0, 16'd20357, 16'd33171, 16'd36685, 16'd47841, 16'd43193, 16'd2465, 16'd59016, 16'd23071, 16'd42671, 16'd57423}; // indx = 3173
    #10;
    addra = 32'd101568;
    dina = {96'd0, 16'd45915, 16'd35986, 16'd21369, 16'd57260, 16'd38630, 16'd17486, 16'd60795, 16'd19138, 16'd30643, 16'd1258}; // indx = 3174
    #10;
    addra = 32'd101600;
    dina = {96'd0, 16'd3488, 16'd3509, 16'd64560, 16'd25991, 16'd1584, 16'd19342, 16'd26743, 16'd9898, 16'd3608, 16'd15768}; // indx = 3175
    #10;
    addra = 32'd101632;
    dina = {96'd0, 16'd20422, 16'd45202, 16'd42395, 16'd57723, 16'd9682, 16'd534, 16'd44226, 16'd14794, 16'd65137, 16'd56181}; // indx = 3176
    #10;
    addra = 32'd101664;
    dina = {96'd0, 16'd23354, 16'd31968, 16'd2483, 16'd28192, 16'd23244, 16'd38835, 16'd45757, 16'd18229, 16'd35454, 16'd32497}; // indx = 3177
    #10;
    addra = 32'd101696;
    dina = {96'd0, 16'd59413, 16'd25580, 16'd33965, 16'd6783, 16'd40908, 16'd54370, 16'd28241, 16'd21217, 16'd9011, 16'd26182}; // indx = 3178
    #10;
    addra = 32'd101728;
    dina = {96'd0, 16'd64735, 16'd15074, 16'd63802, 16'd47295, 16'd23666, 16'd18416, 16'd33912, 16'd39060, 16'd19632, 16'd3147}; // indx = 3179
    #10;
    addra = 32'd101760;
    dina = {96'd0, 16'd8992, 16'd33062, 16'd1025, 16'd51195, 16'd31516, 16'd17277, 16'd42241, 16'd48154, 16'd33668, 16'd48239}; // indx = 3180
    #10;
    addra = 32'd101792;
    dina = {96'd0, 16'd35934, 16'd61331, 16'd38314, 16'd57482, 16'd28388, 16'd26229, 16'd9145, 16'd60149, 16'd13721, 16'd23671}; // indx = 3181
    #10;
    addra = 32'd101824;
    dina = {96'd0, 16'd23432, 16'd29891, 16'd48885, 16'd52563, 16'd20175, 16'd2472, 16'd5660, 16'd9069, 16'd13314, 16'd16975}; // indx = 3182
    #10;
    addra = 32'd101856;
    dina = {96'd0, 16'd640, 16'd42574, 16'd49700, 16'd13852, 16'd56179, 16'd7796, 16'd10485, 16'd51865, 16'd10592, 16'd32025}; // indx = 3183
    #10;
    addra = 32'd101888;
    dina = {96'd0, 16'd57254, 16'd9055, 16'd49404, 16'd63094, 16'd23366, 16'd32150, 16'd37082, 16'd43767, 16'd33562, 16'd41914}; // indx = 3184
    #10;
    addra = 32'd101920;
    dina = {96'd0, 16'd3433, 16'd6531, 16'd27306, 16'd23820, 16'd37592, 16'd40401, 16'd35783, 16'd27493, 16'd24818, 16'd59022}; // indx = 3185
    #10;
    addra = 32'd101952;
    dina = {96'd0, 16'd4720, 16'd58901, 16'd5530, 16'd17798, 16'd6762, 16'd45914, 16'd33266, 16'd2615, 16'd39337, 16'd23920}; // indx = 3186
    #10;
    addra = 32'd101984;
    dina = {96'd0, 16'd52151, 16'd61539, 16'd53293, 16'd19242, 16'd3880, 16'd20977, 16'd64447, 16'd3149, 16'd27212, 16'd26400}; // indx = 3187
    #10;
    addra = 32'd102016;
    dina = {96'd0, 16'd56413, 16'd29677, 16'd13226, 16'd50663, 16'd8819, 16'd9772, 16'd15897, 16'd52671, 16'd20767, 16'd41126}; // indx = 3188
    #10;
    addra = 32'd102048;
    dina = {96'd0, 16'd22655, 16'd6661, 16'd16581, 16'd53982, 16'd6072, 16'd38776, 16'd30459, 16'd61594, 16'd8231, 16'd21686}; // indx = 3189
    #10;
    addra = 32'd102080;
    dina = {96'd0, 16'd46799, 16'd14984, 16'd28955, 16'd64909, 16'd41971, 16'd38795, 16'd25191, 16'd40664, 16'd18776, 16'd14757}; // indx = 3190
    #10;
    addra = 32'd102112;
    dina = {96'd0, 16'd368, 16'd31806, 16'd530, 16'd43841, 16'd43690, 16'd3010, 16'd47809, 16'd60564, 16'd19545, 16'd57264}; // indx = 3191
    #10;
    addra = 32'd102144;
    dina = {96'd0, 16'd4944, 16'd7928, 16'd57014, 16'd2400, 16'd39024, 16'd22093, 16'd44090, 16'd59293, 16'd19918, 16'd43527}; // indx = 3192
    #10;
    addra = 32'd102176;
    dina = {96'd0, 16'd57815, 16'd31518, 16'd60778, 16'd46247, 16'd35238, 16'd42491, 16'd35800, 16'd50077, 16'd10782, 16'd26528}; // indx = 3193
    #10;
    addra = 32'd102208;
    dina = {96'd0, 16'd56336, 16'd37825, 16'd17998, 16'd50564, 16'd33450, 16'd15910, 16'd32928, 16'd28522, 16'd14488, 16'd9152}; // indx = 3194
    #10;
    addra = 32'd102240;
    dina = {96'd0, 16'd39865, 16'd23388, 16'd3183, 16'd28324, 16'd29525, 16'd36880, 16'd17180, 16'd21191, 16'd22721, 16'd51960}; // indx = 3195
    #10;
    addra = 32'd102272;
    dina = {96'd0, 16'd9528, 16'd17661, 16'd61267, 16'd55631, 16'd53112, 16'd34774, 16'd48170, 16'd56757, 16'd23384, 16'd32535}; // indx = 3196
    #10;
    addra = 32'd102304;
    dina = {96'd0, 16'd52148, 16'd5576, 16'd64872, 16'd49922, 16'd19606, 16'd35329, 16'd39178, 16'd56997, 16'd9155, 16'd7987}; // indx = 3197
    #10;
    addra = 32'd102336;
    dina = {96'd0, 16'd36761, 16'd2812, 16'd82, 16'd5328, 16'd38540, 16'd17023, 16'd48942, 16'd4307, 16'd58401, 16'd15334}; // indx = 3198
    #10;
    addra = 32'd102368;
    dina = {96'd0, 16'd53549, 16'd46652, 16'd452, 16'd28512, 16'd8264, 16'd19304, 16'd53674, 16'd11048, 16'd17310, 16'd9136}; // indx = 3199
    #10;
    addra = 32'd102400;
    dina = {96'd0, 16'd40092, 16'd41551, 16'd25217, 16'd55424, 16'd61257, 16'd64904, 16'd19405, 16'd13922, 16'd10748, 16'd48560}; // indx = 3200
    #10;
    addra = 32'd102432;
    dina = {96'd0, 16'd63007, 16'd18161, 16'd15866, 16'd55190, 16'd60293, 16'd34753, 16'd3324, 16'd28870, 16'd43448, 16'd64347}; // indx = 3201
    #10;
    addra = 32'd102464;
    dina = {96'd0, 16'd34708, 16'd54276, 16'd24021, 16'd2058, 16'd5336, 16'd26582, 16'd56934, 16'd52887, 16'd50460, 16'd30789}; // indx = 3202
    #10;
    addra = 32'd102496;
    dina = {96'd0, 16'd51086, 16'd30453, 16'd24607, 16'd37456, 16'd56510, 16'd65271, 16'd6544, 16'd24112, 16'd9665, 16'd4266}; // indx = 3203
    #10;
    addra = 32'd102528;
    dina = {96'd0, 16'd18211, 16'd4013, 16'd59324, 16'd1365, 16'd57959, 16'd23405, 16'd36515, 16'd5405, 16'd22161, 16'd32385}; // indx = 3204
    #10;
    addra = 32'd102560;
    dina = {96'd0, 16'd47630, 16'd34849, 16'd39448, 16'd35166, 16'd64031, 16'd1875, 16'd37368, 16'd48700, 16'd47476, 16'd41981}; // indx = 3205
    #10;
    addra = 32'd102592;
    dina = {96'd0, 16'd46658, 16'd32367, 16'd24083, 16'd27942, 16'd16241, 16'd15287, 16'd15748, 16'd1982, 16'd19938, 16'd53525}; // indx = 3206
    #10;
    addra = 32'd102624;
    dina = {96'd0, 16'd57144, 16'd12304, 16'd34607, 16'd49963, 16'd22195, 16'd46844, 16'd22987, 16'd39112, 16'd43175, 16'd55764}; // indx = 3207
    #10;
    addra = 32'd102656;
    dina = {96'd0, 16'd23840, 16'd31644, 16'd34356, 16'd56560, 16'd1460, 16'd3245, 16'd868, 16'd63310, 16'd48977, 16'd42160}; // indx = 3208
    #10;
    addra = 32'd102688;
    dina = {96'd0, 16'd13151, 16'd54511, 16'd3252, 16'd42581, 16'd39330, 16'd4968, 16'd60969, 16'd24367, 16'd56541, 16'd27762}; // indx = 3209
    #10;
    addra = 32'd102720;
    dina = {96'd0, 16'd31450, 16'd46944, 16'd13836, 16'd47300, 16'd47136, 16'd8840, 16'd37015, 16'd60271, 16'd20193, 16'd27755}; // indx = 3210
    #10;
    addra = 32'd102752;
    dina = {96'd0, 16'd38592, 16'd63599, 16'd254, 16'd20809, 16'd9209, 16'd15001, 16'd56266, 16'd24358, 16'd36085, 16'd31234}; // indx = 3211
    #10;
    addra = 32'd102784;
    dina = {96'd0, 16'd24715, 16'd13847, 16'd49611, 16'd35926, 16'd64920, 16'd45803, 16'd55622, 16'd49340, 16'd3076, 16'd2722}; // indx = 3212
    #10;
    addra = 32'd102816;
    dina = {96'd0, 16'd5064, 16'd18728, 16'd12621, 16'd17906, 16'd55158, 16'd30522, 16'd4474, 16'd3815, 16'd49656, 16'd62657}; // indx = 3213
    #10;
    addra = 32'd102848;
    dina = {96'd0, 16'd9170, 16'd12107, 16'd15269, 16'd12434, 16'd61256, 16'd46061, 16'd27318, 16'd6716, 16'd5779, 16'd17577}; // indx = 3214
    #10;
    addra = 32'd102880;
    dina = {96'd0, 16'd39648, 16'd58346, 16'd19341, 16'd55942, 16'd20607, 16'd24484, 16'd35622, 16'd33472, 16'd22588, 16'd34600}; // indx = 3215
    #10;
    addra = 32'd102912;
    dina = {96'd0, 16'd21482, 16'd28170, 16'd40188, 16'd17859, 16'd43163, 16'd26242, 16'd27658, 16'd10498, 16'd35144, 16'd25127}; // indx = 3216
    #10;
    addra = 32'd102944;
    dina = {96'd0, 16'd15282, 16'd52095, 16'd55307, 16'd38622, 16'd45606, 16'd55784, 16'd38932, 16'd11288, 16'd22221, 16'd12785}; // indx = 3217
    #10;
    addra = 32'd102976;
    dina = {96'd0, 16'd6768, 16'd41307, 16'd14914, 16'd52537, 16'd28788, 16'd39036, 16'd1510, 16'd61320, 16'd21096, 16'd4460}; // indx = 3218
    #10;
    addra = 32'd103008;
    dina = {96'd0, 16'd25810, 16'd24849, 16'd55405, 16'd30083, 16'd38555, 16'd11351, 16'd58988, 16'd28339, 16'd15494, 16'd25067}; // indx = 3219
    #10;
    addra = 32'd103040;
    dina = {96'd0, 16'd60634, 16'd20389, 16'd9010, 16'd12788, 16'd39757, 16'd63588, 16'd11346, 16'd64469, 16'd50502, 16'd17733}; // indx = 3220
    #10;
    addra = 32'd103072;
    dina = {96'd0, 16'd18022, 16'd6230, 16'd958, 16'd53998, 16'd2989, 16'd16321, 16'd32485, 16'd4050, 16'd21488, 16'd36675}; // indx = 3221
    #10;
    addra = 32'd103104;
    dina = {96'd0, 16'd19012, 16'd20485, 16'd145, 16'd44279, 16'd16181, 16'd26399, 16'd40238, 16'd40171, 16'd59498, 16'd45079}; // indx = 3222
    #10;
    addra = 32'd103136;
    dina = {96'd0, 16'd39042, 16'd51035, 16'd15199, 16'd5617, 16'd278, 16'd5208, 16'd63406, 16'd43314, 16'd42686, 16'd13110}; // indx = 3223
    #10;
    addra = 32'd103168;
    dina = {96'd0, 16'd60881, 16'd44792, 16'd30524, 16'd19286, 16'd47334, 16'd20670, 16'd33809, 16'd8084, 16'd28415, 16'd9790}; // indx = 3224
    #10;
    addra = 32'd103200;
    dina = {96'd0, 16'd21426, 16'd1667, 16'd9831, 16'd55772, 16'd19654, 16'd54581, 16'd24831, 16'd13945, 16'd40764, 16'd11022}; // indx = 3225
    #10;
    addra = 32'd103232;
    dina = {96'd0, 16'd34281, 16'd10915, 16'd59274, 16'd21209, 16'd39883, 16'd17036, 16'd62830, 16'd12067, 16'd10670, 16'd15082}; // indx = 3226
    #10;
    addra = 32'd103264;
    dina = {96'd0, 16'd34712, 16'd384, 16'd46421, 16'd45433, 16'd33801, 16'd31716, 16'd64067, 16'd57293, 16'd40617, 16'd1389}; // indx = 3227
    #10;
    addra = 32'd103296;
    dina = {96'd0, 16'd43062, 16'd21542, 16'd48112, 16'd4359, 16'd17610, 16'd4596, 16'd25540, 16'd37315, 16'd53639, 16'd43821}; // indx = 3228
    #10;
    addra = 32'd103328;
    dina = {96'd0, 16'd26927, 16'd48744, 16'd61775, 16'd48663, 16'd17198, 16'd4515, 16'd44309, 16'd63620, 16'd14563, 16'd51326}; // indx = 3229
    #10;
    addra = 32'd103360;
    dina = {96'd0, 16'd27081, 16'd37451, 16'd50882, 16'd25985, 16'd48791, 16'd48956, 16'd17938, 16'd47416, 16'd57568, 16'd20174}; // indx = 3230
    #10;
    addra = 32'd103392;
    dina = {96'd0, 16'd1026, 16'd9237, 16'd15022, 16'd2400, 16'd22640, 16'd54931, 16'd59265, 16'd26774, 16'd44830, 16'd20747}; // indx = 3231
    #10;
    addra = 32'd103424;
    dina = {96'd0, 16'd9156, 16'd2809, 16'd13516, 16'd17121, 16'd9508, 16'd51489, 16'd1301, 16'd25113, 16'd7635, 16'd53995}; // indx = 3232
    #10;
    addra = 32'd103456;
    dina = {96'd0, 16'd53554, 16'd44816, 16'd56756, 16'd15579, 16'd51662, 16'd12862, 16'd45834, 16'd23973, 16'd54056, 16'd57881}; // indx = 3233
    #10;
    addra = 32'd103488;
    dina = {96'd0, 16'd65182, 16'd19036, 16'd20829, 16'd40064, 16'd37928, 16'd9571, 16'd31983, 16'd41581, 16'd26683, 16'd26131}; // indx = 3234
    #10;
    addra = 32'd103520;
    dina = {96'd0, 16'd46866, 16'd42347, 16'd1015, 16'd11903, 16'd57086, 16'd57586, 16'd13089, 16'd16180, 16'd17879, 16'd34683}; // indx = 3235
    #10;
    addra = 32'd103552;
    dina = {96'd0, 16'd50103, 16'd55453, 16'd7637, 16'd26460, 16'd1272, 16'd57025, 16'd14915, 16'd42817, 16'd56793, 16'd20424}; // indx = 3236
    #10;
    addra = 32'd103584;
    dina = {96'd0, 16'd47748, 16'd36067, 16'd1824, 16'd15016, 16'd34967, 16'd36701, 16'd40114, 16'd51784, 16'd41977, 16'd58468}; // indx = 3237
    #10;
    addra = 32'd103616;
    dina = {96'd0, 16'd56968, 16'd23846, 16'd12742, 16'd34465, 16'd22092, 16'd13292, 16'd20180, 16'd31277, 16'd59702, 16'd7008}; // indx = 3238
    #10;
    addra = 32'd103648;
    dina = {96'd0, 16'd12775, 16'd50910, 16'd51530, 16'd12539, 16'd7580, 16'd15004, 16'd44308, 16'd42900, 16'd3212, 16'd62400}; // indx = 3239
    #10;
    addra = 32'd103680;
    dina = {96'd0, 16'd58186, 16'd42017, 16'd56480, 16'd1562, 16'd13480, 16'd9088, 16'd53861, 16'd3130, 16'd12383, 16'd19703}; // indx = 3240
    #10;
    addra = 32'd103712;
    dina = {96'd0, 16'd59852, 16'd51762, 16'd28845, 16'd50999, 16'd5864, 16'd29005, 16'd23819, 16'd3175, 16'd34269, 16'd12265}; // indx = 3241
    #10;
    addra = 32'd103744;
    dina = {96'd0, 16'd40213, 16'd46381, 16'd29128, 16'd28565, 16'd20089, 16'd17895, 16'd12091, 16'd45068, 16'd57647, 16'd37291}; // indx = 3242
    #10;
    addra = 32'd103776;
    dina = {96'd0, 16'd48619, 16'd46994, 16'd44780, 16'd58070, 16'd8510, 16'd12319, 16'd50035, 16'd5916, 16'd14241, 16'd19305}; // indx = 3243
    #10;
    addra = 32'd103808;
    dina = {96'd0, 16'd36841, 16'd62089, 16'd64284, 16'd62871, 16'd46033, 16'd22674, 16'd60251, 16'd19563, 16'd43359, 16'd31110}; // indx = 3244
    #10;
    addra = 32'd103840;
    dina = {96'd0, 16'd54480, 16'd6532, 16'd59809, 16'd5544, 16'd1262, 16'd24110, 16'd2607, 16'd42701, 16'd23772, 16'd21067}; // indx = 3245
    #10;
    addra = 32'd103872;
    dina = {96'd0, 16'd45811, 16'd3368, 16'd1515, 16'd31103, 16'd40911, 16'd10381, 16'd892, 16'd53180, 16'd15072, 16'd17569}; // indx = 3246
    #10;
    addra = 32'd103904;
    dina = {96'd0, 16'd7400, 16'd38313, 16'd6923, 16'd37453, 16'd886, 16'd7192, 16'd32192, 16'd12827, 16'd53874, 16'd19075}; // indx = 3247
    #10;
    addra = 32'd103936;
    dina = {96'd0, 16'd55435, 16'd56682, 16'd48210, 16'd49997, 16'd45999, 16'd5621, 16'd45345, 16'd53071, 16'd26018, 16'd5827}; // indx = 3248
    #10;
    addra = 32'd103968;
    dina = {96'd0, 16'd27629, 16'd24434, 16'd54661, 16'd7051, 16'd52412, 16'd61657, 16'd8198, 16'd21345, 16'd42251, 16'd55435}; // indx = 3249
    #10;
    addra = 32'd104000;
    dina = {96'd0, 16'd52285, 16'd28767, 16'd48406, 16'd57555, 16'd42053, 16'd12301, 16'd60590, 16'd19570, 16'd4295, 16'd55405}; // indx = 3250
    #10;
    addra = 32'd104032;
    dina = {96'd0, 16'd27477, 16'd60275, 16'd9527, 16'd35443, 16'd1327, 16'd60070, 16'd58299, 16'd64746, 16'd44949, 16'd42037}; // indx = 3251
    #10;
    addra = 32'd104064;
    dina = {96'd0, 16'd55336, 16'd45076, 16'd54660, 16'd1742, 16'd34342, 16'd43972, 16'd40529, 16'd49349, 16'd12012, 16'd64286}; // indx = 3252
    #10;
    addra = 32'd104096;
    dina = {96'd0, 16'd32049, 16'd24653, 16'd7480, 16'd32908, 16'd3568, 16'd46372, 16'd43218, 16'd31093, 16'd61130, 16'd46713}; // indx = 3253
    #10;
    addra = 32'd104128;
    dina = {96'd0, 16'd38229, 16'd15490, 16'd38502, 16'd52638, 16'd1511, 16'd62058, 16'd27369, 16'd13986, 16'd4416, 16'd53211}; // indx = 3254
    #10;
    addra = 32'd104160;
    dina = {96'd0, 16'd28880, 16'd47648, 16'd55440, 16'd50122, 16'd60343, 16'd9399, 16'd15401, 16'd24096, 16'd10414, 16'd26502}; // indx = 3255
    #10;
    addra = 32'd104192;
    dina = {96'd0, 16'd18575, 16'd25065, 16'd11923, 16'd21110, 16'd40839, 16'd28178, 16'd37005, 16'd10566, 16'd29912, 16'd25838}; // indx = 3256
    #10;
    addra = 32'd104224;
    dina = {96'd0, 16'd54945, 16'd42538, 16'd54287, 16'd16240, 16'd51821, 16'd5735, 16'd21355, 16'd29366, 16'd64731, 16'd4906}; // indx = 3257
    #10;
    addra = 32'd104256;
    dina = {96'd0, 16'd24881, 16'd28128, 16'd30232, 16'd55288, 16'd13206, 16'd44312, 16'd55378, 16'd4298, 16'd12236, 16'd49867}; // indx = 3258
    #10;
    addra = 32'd104288;
    dina = {96'd0, 16'd12644, 16'd58558, 16'd11184, 16'd50190, 16'd4553, 16'd8690, 16'd41412, 16'd39994, 16'd53169, 16'd38587}; // indx = 3259
    #10;
    addra = 32'd104320;
    dina = {96'd0, 16'd15521, 16'd20558, 16'd52639, 16'd2481, 16'd55623, 16'd28566, 16'd53328, 16'd18101, 16'd21748, 16'd26163}; // indx = 3260
    #10;
    addra = 32'd104352;
    dina = {96'd0, 16'd49196, 16'd12992, 16'd50280, 16'd9753, 16'd1115, 16'd3129, 16'd64084, 16'd409, 16'd1208, 16'd61426}; // indx = 3261
    #10;
    addra = 32'd104384;
    dina = {96'd0, 16'd64744, 16'd30344, 16'd27184, 16'd26348, 16'd35539, 16'd60752, 16'd12425, 16'd46082, 16'd7263, 16'd4446}; // indx = 3262
    #10;
    addra = 32'd104416;
    dina = {96'd0, 16'd16715, 16'd21638, 16'd57532, 16'd29384, 16'd28464, 16'd14953, 16'd13762, 16'd37398, 16'd7885, 16'd50440}; // indx = 3263
    #10;
    addra = 32'd104448;
    dina = {96'd0, 16'd20093, 16'd52709, 16'd48585, 16'd62199, 16'd52926, 16'd43825, 16'd14582, 16'd37143, 16'd38421, 16'd59588}; // indx = 3264
    #10;
    addra = 32'd104480;
    dina = {96'd0, 16'd39365, 16'd5853, 16'd62351, 16'd47006, 16'd20059, 16'd21843, 16'd9662, 16'd24749, 16'd4137, 16'd36129}; // indx = 3265
    #10;
    addra = 32'd104512;
    dina = {96'd0, 16'd1244, 16'd29234, 16'd12868, 16'd39672, 16'd48727, 16'd12263, 16'd9272, 16'd10064, 16'd36970, 16'd56709}; // indx = 3266
    #10;
    addra = 32'd104544;
    dina = {96'd0, 16'd4464, 16'd35521, 16'd4907, 16'd56302, 16'd62814, 16'd59051, 16'd41608, 16'd48124, 16'd39129, 16'd52074}; // indx = 3267
    #10;
    addra = 32'd104576;
    dina = {96'd0, 16'd19733, 16'd34036, 16'd57776, 16'd46803, 16'd53117, 16'd2513, 16'd47355, 16'd10335, 16'd44822, 16'd39510}; // indx = 3268
    #10;
    addra = 32'd104608;
    dina = {96'd0, 16'd53824, 16'd18781, 16'd49442, 16'd45649, 16'd18875, 16'd266, 16'd50624, 16'd41253, 16'd4270, 16'd47036}; // indx = 3269
    #10;
    addra = 32'd104640;
    dina = {96'd0, 16'd44792, 16'd58914, 16'd2831, 16'd6288, 16'd23834, 16'd48375, 16'd51262, 16'd49271, 16'd40699, 16'd32534}; // indx = 3270
    #10;
    addra = 32'd104672;
    dina = {96'd0, 16'd46137, 16'd32584, 16'd38862, 16'd45499, 16'd25408, 16'd18101, 16'd3514, 16'd62402, 16'd36468, 16'd21055}; // indx = 3271
    #10;
    addra = 32'd104704;
    dina = {96'd0, 16'd2785, 16'd55977, 16'd50757, 16'd42415, 16'd16478, 16'd28200, 16'd11463, 16'd35083, 16'd1623, 16'd52387}; // indx = 3272
    #10;
    addra = 32'd104736;
    dina = {96'd0, 16'd6593, 16'd45874, 16'd42496, 16'd49325, 16'd19128, 16'd13555, 16'd18155, 16'd37262, 16'd23113, 16'd2997}; // indx = 3273
    #10;
    addra = 32'd104768;
    dina = {96'd0, 16'd48850, 16'd42944, 16'd18771, 16'd41379, 16'd33586, 16'd22748, 16'd26105, 16'd62131, 16'd15641, 16'd10769}; // indx = 3274
    #10;
    addra = 32'd104800;
    dina = {96'd0, 16'd41046, 16'd13853, 16'd17560, 16'd48832, 16'd3262, 16'd42936, 16'd51288, 16'd63546, 16'd3507, 16'd40034}; // indx = 3275
    #10;
    addra = 32'd104832;
    dina = {96'd0, 16'd54636, 16'd28865, 16'd10494, 16'd9155, 16'd34552, 16'd64381, 16'd3874, 16'd45496, 16'd55051, 16'd45798}; // indx = 3276
    #10;
    addra = 32'd104864;
    dina = {96'd0, 16'd52729, 16'd12638, 16'd13867, 16'd46025, 16'd12187, 16'd996, 16'd53060, 16'd16784, 16'd36737, 16'd51323}; // indx = 3277
    #10;
    addra = 32'd104896;
    dina = {96'd0, 16'd36500, 16'd17978, 16'd57163, 16'd22273, 16'd45706, 16'd4082, 16'd20729, 16'd30875, 16'd59751, 16'd40461}; // indx = 3278
    #10;
    addra = 32'd104928;
    dina = {96'd0, 16'd63320, 16'd42019, 16'd59612, 16'd60499, 16'd58262, 16'd9888, 16'd11947, 16'd2707, 16'd43855, 16'd29924}; // indx = 3279
    #10;
    addra = 32'd104960;
    dina = {96'd0, 16'd18448, 16'd38623, 16'd50951, 16'd5715, 16'd59164, 16'd50378, 16'd44428, 16'd31884, 16'd25957, 16'd35129}; // indx = 3280
    #10;
    addra = 32'd104992;
    dina = {96'd0, 16'd47832, 16'd11952, 16'd34311, 16'd38681, 16'd7046, 16'd30062, 16'd60621, 16'd42115, 16'd27987, 16'd51773}; // indx = 3281
    #10;
    addra = 32'd105024;
    dina = {96'd0, 16'd54881, 16'd8326, 16'd57091, 16'd9028, 16'd64464, 16'd8122, 16'd32363, 16'd35985, 16'd21266, 16'd61660}; // indx = 3282
    #10;
    addra = 32'd105056;
    dina = {96'd0, 16'd21200, 16'd8252, 16'd4015, 16'd16633, 16'd58822, 16'd56675, 16'd32501, 16'd15546, 16'd28743, 16'd55653}; // indx = 3283
    #10;
    addra = 32'd105088;
    dina = {96'd0, 16'd55151, 16'd56560, 16'd51604, 16'd54584, 16'd31943, 16'd28967, 16'd13782, 16'd40805, 16'd57414, 16'd24330}; // indx = 3284
    #10;
    addra = 32'd105120;
    dina = {96'd0, 16'd10414, 16'd15164, 16'd59028, 16'd12884, 16'd22512, 16'd58813, 16'd26663, 16'd12792, 16'd8357, 16'd33937}; // indx = 3285
    #10;
    addra = 32'd105152;
    dina = {96'd0, 16'd49850, 16'd43751, 16'd57200, 16'd33157, 16'd10002, 16'd25130, 16'd18010, 16'd599, 16'd29460, 16'd19774}; // indx = 3286
    #10;
    addra = 32'd105184;
    dina = {96'd0, 16'd18547, 16'd7854, 16'd19067, 16'd53691, 16'd29514, 16'd37591, 16'd63176, 16'd43052, 16'd2166, 16'd36168}; // indx = 3287
    #10;
    addra = 32'd105216;
    dina = {96'd0, 16'd13617, 16'd60251, 16'd35599, 16'd35325, 16'd60561, 16'd26053, 16'd52802, 16'd53785, 16'd6266, 16'd43547}; // indx = 3288
    #10;
    addra = 32'd105248;
    dina = {96'd0, 16'd13513, 16'd9282, 16'd15216, 16'd37677, 16'd59005, 16'd51172, 16'd28575, 16'd59052, 16'd54194, 16'd19196}; // indx = 3289
    #10;
    addra = 32'd105280;
    dina = {96'd0, 16'd33379, 16'd24500, 16'd14905, 16'd8034, 16'd33828, 16'd757, 16'd54607, 16'd32011, 16'd16761, 16'd60386}; // indx = 3290
    #10;
    addra = 32'd105312;
    dina = {96'd0, 16'd52169, 16'd48728, 16'd19080, 16'd24160, 16'd41472, 16'd24667, 16'd41118, 16'd19375, 16'd21354, 16'd48277}; // indx = 3291
    #10;
    addra = 32'd105344;
    dina = {96'd0, 16'd33150, 16'd22358, 16'd47223, 16'd28857, 16'd13703, 16'd58355, 16'd20961, 16'd15358, 16'd45681, 16'd16980}; // indx = 3292
    #10;
    addra = 32'd105376;
    dina = {96'd0, 16'd27755, 16'd49220, 16'd9097, 16'd30228, 16'd23421, 16'd41477, 16'd37874, 16'd27781, 16'd30024, 16'd55281}; // indx = 3293
    #10;
    addra = 32'd105408;
    dina = {96'd0, 16'd41081, 16'd24489, 16'd54214, 16'd5194, 16'd39732, 16'd58376, 16'd56053, 16'd32629, 16'd5245, 16'd39113}; // indx = 3294
    #10;
    addra = 32'd105440;
    dina = {96'd0, 16'd46422, 16'd32632, 16'd16916, 16'd58807, 16'd1513, 16'd21781, 16'd21699, 16'd16295, 16'd3319, 16'd26138}; // indx = 3295
    #10;
    addra = 32'd105472;
    dina = {96'd0, 16'd38786, 16'd37669, 16'd9570, 16'd49053, 16'd30337, 16'd65284, 16'd31455, 16'd64807, 16'd49744, 16'd58902}; // indx = 3296
    #10;
    addra = 32'd105504;
    dina = {96'd0, 16'd50594, 16'd9713, 16'd15934, 16'd33697, 16'd36433, 16'd17315, 16'd28621, 16'd25795, 16'd33164, 16'd28450}; // indx = 3297
    #10;
    addra = 32'd105536;
    dina = {96'd0, 16'd49839, 16'd40417, 16'd36080, 16'd28243, 16'd13592, 16'd5237, 16'd19084, 16'd38445, 16'd58228, 16'd37185}; // indx = 3298
    #10;
    addra = 32'd105568;
    dina = {96'd0, 16'd49775, 16'd48707, 16'd29654, 16'd24723, 16'd59920, 16'd21012, 16'd25234, 16'd11095, 16'd37155, 16'd30015}; // indx = 3299
    #10;
    addra = 32'd105600;
    dina = {96'd0, 16'd57844, 16'd65030, 16'd31625, 16'd12676, 16'd415, 16'd48820, 16'd57492, 16'd55669, 16'd38758, 16'd47042}; // indx = 3300
    #10;
    addra = 32'd105632;
    dina = {96'd0, 16'd219, 16'd65280, 16'd38607, 16'd62508, 16'd65343, 16'd12516, 16'd46006, 16'd17844, 16'd15519, 16'd22993}; // indx = 3301
    #10;
    addra = 32'd105664;
    dina = {96'd0, 16'd18896, 16'd61644, 16'd29114, 16'd19187, 16'd50111, 16'd2553, 16'd39686, 16'd20733, 16'd5821, 16'd7447}; // indx = 3302
    #10;
    addra = 32'd105696;
    dina = {96'd0, 16'd1170, 16'd33414, 16'd16954, 16'd44865, 16'd63489, 16'd22404, 16'd22001, 16'd29543, 16'd63050, 16'd50333}; // indx = 3303
    #10;
    addra = 32'd105728;
    dina = {96'd0, 16'd12461, 16'd10563, 16'd1796, 16'd29430, 16'd26605, 16'd34805, 16'd38063, 16'd25884, 16'd5409, 16'd41385}; // indx = 3304
    #10;
    addra = 32'd105760;
    dina = {96'd0, 16'd25492, 16'd31446, 16'd802, 16'd11561, 16'd24576, 16'd25111, 16'd33556, 16'd17147, 16'd55280, 16'd5626}; // indx = 3305
    #10;
    addra = 32'd105792;
    dina = {96'd0, 16'd4222, 16'd54879, 16'd49083, 16'd31439, 16'd26403, 16'd63340, 16'd47619, 16'd61516, 16'd16495, 16'd42477}; // indx = 3306
    #10;
    addra = 32'd105824;
    dina = {96'd0, 16'd51517, 16'd29610, 16'd2258, 16'd1037, 16'd2605, 16'd40140, 16'd14010, 16'd64286, 16'd36616, 16'd61268}; // indx = 3307
    #10;
    addra = 32'd105856;
    dina = {96'd0, 16'd4111, 16'd49189, 16'd47401, 16'd50250, 16'd58383, 16'd48618, 16'd27745, 16'd41006, 16'd25927, 16'd63106}; // indx = 3308
    #10;
    addra = 32'd105888;
    dina = {96'd0, 16'd24893, 16'd20597, 16'd29271, 16'd44625, 16'd43950, 16'd53024, 16'd36577, 16'd34132, 16'd63900, 16'd51927}; // indx = 3309
    #10;
    addra = 32'd105920;
    dina = {96'd0, 16'd61163, 16'd35234, 16'd64170, 16'd64515, 16'd9597, 16'd56779, 16'd42339, 16'd6142, 16'd54319, 16'd8513}; // indx = 3310
    #10;
    addra = 32'd105952;
    dina = {96'd0, 16'd21220, 16'd29401, 16'd49225, 16'd31148, 16'd1057, 16'd7387, 16'd48945, 16'd58780, 16'd53522, 16'd25184}; // indx = 3311
    #10;
    addra = 32'd105984;
    dina = {96'd0, 16'd5825, 16'd20018, 16'd49899, 16'd24689, 16'd14186, 16'd40407, 16'd19936, 16'd61755, 16'd27192, 16'd59869}; // indx = 3312
    #10;
    addra = 32'd106016;
    dina = {96'd0, 16'd59429, 16'd6521, 16'd4261, 16'd49996, 16'd17805, 16'd12258, 16'd49526, 16'd45482, 16'd5354, 16'd64404}; // indx = 3313
    #10;
    addra = 32'd106048;
    dina = {96'd0, 16'd828, 16'd54051, 16'd56853, 16'd21818, 16'd32900, 16'd11350, 16'd62412, 16'd32439, 16'd54377, 16'd23202}; // indx = 3314
    #10;
    addra = 32'd106080;
    dina = {96'd0, 16'd18762, 16'd45343, 16'd61003, 16'd30609, 16'd55855, 16'd36631, 16'd18061, 16'd54759, 16'd24955, 16'd31261}; // indx = 3315
    #10;
    addra = 32'd106112;
    dina = {96'd0, 16'd18696, 16'd44636, 16'd13207, 16'd9516, 16'd35063, 16'd37471, 16'd40305, 16'd33642, 16'd1488, 16'd41205}; // indx = 3316
    #10;
    addra = 32'd106144;
    dina = {96'd0, 16'd45461, 16'd61386, 16'd61486, 16'd34684, 16'd33694, 16'd40026, 16'd45852, 16'd18020, 16'd39726, 16'd19347}; // indx = 3317
    #10;
    addra = 32'd106176;
    dina = {96'd0, 16'd15586, 16'd52667, 16'd1502, 16'd54545, 16'd63757, 16'd40681, 16'd4155, 16'd51621, 16'd27184, 16'd45305}; // indx = 3318
    #10;
    addra = 32'd106208;
    dina = {96'd0, 16'd47469, 16'd63640, 16'd53857, 16'd25115, 16'd6632, 16'd59839, 16'd10099, 16'd9622, 16'd23584, 16'd38846}; // indx = 3319
    #10;
    addra = 32'd106240;
    dina = {96'd0, 16'd54885, 16'd3667, 16'd59309, 16'd50057, 16'd59164, 16'd45469, 16'd5045, 16'd36730, 16'd42870, 16'd64158}; // indx = 3320
    #10;
    addra = 32'd106272;
    dina = {96'd0, 16'd26660, 16'd44442, 16'd49468, 16'd37795, 16'd40477, 16'd9685, 16'd58053, 16'd10818, 16'd46879, 16'd37846}; // indx = 3321
    #10;
    addra = 32'd106304;
    dina = {96'd0, 16'd5735, 16'd36705, 16'd21616, 16'd56944, 16'd36391, 16'd29269, 16'd38091, 16'd25848, 16'd55326, 16'd46513}; // indx = 3322
    #10;
    addra = 32'd106336;
    dina = {96'd0, 16'd55205, 16'd40274, 16'd51940, 16'd43417, 16'd5200, 16'd41838, 16'd3801, 16'd52064, 16'd37022, 16'd12587}; // indx = 3323
    #10;
    addra = 32'd106368;
    dina = {96'd0, 16'd63190, 16'd27935, 16'd10581, 16'd11574, 16'd57306, 16'd46480, 16'd64800, 16'd63214, 16'd47411, 16'd35193}; // indx = 3324
    #10;
    addra = 32'd106400;
    dina = {96'd0, 16'd48321, 16'd10355, 16'd26280, 16'd46572, 16'd62984, 16'd34998, 16'd48655, 16'd6469, 16'd15203, 16'd46416}; // indx = 3325
    #10;
    addra = 32'd106432;
    dina = {96'd0, 16'd57036, 16'd30433, 16'd35589, 16'd46916, 16'd49235, 16'd1932, 16'd57651, 16'd28054, 16'd24176, 16'd33293}; // indx = 3326
    #10;
    addra = 32'd106464;
    dina = {96'd0, 16'd28184, 16'd24069, 16'd35642, 16'd35853, 16'd55162, 16'd19015, 16'd29813, 16'd52012, 16'd19622, 16'd12944}; // indx = 3327
    #10;
    addra = 32'd106496;
    dina = {96'd0, 16'd53788, 16'd10476, 16'd19253, 16'd62989, 16'd62773, 16'd19352, 16'd19560, 16'd29315, 16'd25105, 16'd55183}; // indx = 3328
    #10;
    addra = 32'd106528;
    dina = {96'd0, 16'd29979, 16'd15243, 16'd39178, 16'd40850, 16'd34405, 16'd13479, 16'd25768, 16'd33704, 16'd31509, 16'd11723}; // indx = 3329
    #10;
    addra = 32'd106560;
    dina = {96'd0, 16'd41298, 16'd47539, 16'd45271, 16'd54744, 16'd49101, 16'd2065, 16'd10243, 16'd28677, 16'd57324, 16'd65173}; // indx = 3330
    #10;
    addra = 32'd106592;
    dina = {96'd0, 16'd55395, 16'd1568, 16'd2941, 16'd47265, 16'd8248, 16'd48964, 16'd6068, 16'd16297, 16'd25039, 16'd22597}; // indx = 3331
    #10;
    addra = 32'd106624;
    dina = {96'd0, 16'd23338, 16'd28810, 16'd45611, 16'd55643, 16'd1309, 16'd41761, 16'd55331, 16'd10454, 16'd22137, 16'd22847}; // indx = 3332
    #10;
    addra = 32'd106656;
    dina = {96'd0, 16'd3009, 16'd35397, 16'd18417, 16'd36567, 16'd14598, 16'd16929, 16'd34413, 16'd11817, 16'd32060, 16'd1987}; // indx = 3333
    #10;
    addra = 32'd106688;
    dina = {96'd0, 16'd32462, 16'd36672, 16'd17796, 16'd43331, 16'd8905, 16'd43278, 16'd12723, 16'd56220, 16'd47331, 16'd19249}; // indx = 3334
    #10;
    addra = 32'd106720;
    dina = {96'd0, 16'd231, 16'd1169, 16'd17139, 16'd52080, 16'd41804, 16'd47308, 16'd16921, 16'd55893, 16'd15844, 16'd46748}; // indx = 3335
    #10;
    addra = 32'd106752;
    dina = {96'd0, 16'd29288, 16'd38039, 16'd12647, 16'd17007, 16'd26487, 16'd1507, 16'd25499, 16'd59581, 16'd20042, 16'd7083}; // indx = 3336
    #10;
    addra = 32'd106784;
    dina = {96'd0, 16'd33718, 16'd23100, 16'd33412, 16'd44062, 16'd32819, 16'd59646, 16'd9130, 16'd53638, 16'd12509, 16'd21330}; // indx = 3337
    #10;
    addra = 32'd106816;
    dina = {96'd0, 16'd37590, 16'd13424, 16'd45165, 16'd54987, 16'd42032, 16'd51414, 16'd10192, 16'd44038, 16'd14219, 16'd21068}; // indx = 3338
    #10;
    addra = 32'd106848;
    dina = {96'd0, 16'd20563, 16'd2665, 16'd36632, 16'd61165, 16'd9198, 16'd30910, 16'd20450, 16'd18252, 16'd37076, 16'd37377}; // indx = 3339
    #10;
    addra = 32'd106880;
    dina = {96'd0, 16'd56102, 16'd30474, 16'd29239, 16'd42799, 16'd40338, 16'd49803, 16'd47983, 16'd37104, 16'd57163, 16'd52056}; // indx = 3340
    #10;
    addra = 32'd106912;
    dina = {96'd0, 16'd49730, 16'd53499, 16'd33788, 16'd53933, 16'd64642, 16'd55496, 16'd55548, 16'd40156, 16'd20576, 16'd59706}; // indx = 3341
    #10;
    addra = 32'd106944;
    dina = {96'd0, 16'd34548, 16'd28800, 16'd16425, 16'd62655, 16'd53400, 16'd45369, 16'd33998, 16'd39269, 16'd38807, 16'd35970}; // indx = 3342
    #10;
    addra = 32'd106976;
    dina = {96'd0, 16'd26809, 16'd22678, 16'd48380, 16'd17991, 16'd62004, 16'd31430, 16'd60859, 16'd63908, 16'd15663, 16'd19210}; // indx = 3343
    #10;
    addra = 32'd107008;
    dina = {96'd0, 16'd44871, 16'd6268, 16'd28098, 16'd4182, 16'd8825, 16'd19957, 16'd33593, 16'd11381, 16'd43560, 16'd30739}; // indx = 3344
    #10;
    addra = 32'd107040;
    dina = {96'd0, 16'd35880, 16'd33015, 16'd12035, 16'd767, 16'd30282, 16'd61125, 16'd17853, 16'd65284, 16'd10915, 16'd25518}; // indx = 3345
    #10;
    addra = 32'd107072;
    dina = {96'd0, 16'd21103, 16'd19496, 16'd5236, 16'd18966, 16'd34985, 16'd50052, 16'd45222, 16'd48936, 16'd48941, 16'd18285}; // indx = 3346
    #10;
    addra = 32'd107104;
    dina = {96'd0, 16'd63378, 16'd22639, 16'd50258, 16'd5082, 16'd45688, 16'd34729, 16'd39124, 16'd22034, 16'd33625, 16'd54998}; // indx = 3347
    #10;
    addra = 32'd107136;
    dina = {96'd0, 16'd29404, 16'd24402, 16'd40088, 16'd5563, 16'd7657, 16'd34026, 16'd16302, 16'd59562, 16'd51965, 16'd40333}; // indx = 3348
    #10;
    addra = 32'd107168;
    dina = {96'd0, 16'd41624, 16'd28985, 16'd50479, 16'd27795, 16'd54424, 16'd39017, 16'd62811, 16'd58903, 16'd56878, 16'd63748}; // indx = 3349
    #10;
    addra = 32'd107200;
    dina = {96'd0, 16'd10877, 16'd21090, 16'd36830, 16'd615, 16'd5164, 16'd31322, 16'd65107, 16'd56072, 16'd27904, 16'd60840}; // indx = 3350
    #10;
    addra = 32'd107232;
    dina = {96'd0, 16'd55485, 16'd16011, 16'd48930, 16'd54793, 16'd7529, 16'd32839, 16'd13008, 16'd13982, 16'd63337, 16'd1401}; // indx = 3351
    #10;
    addra = 32'd107264;
    dina = {96'd0, 16'd2381, 16'd59682, 16'd11762, 16'd28049, 16'd16911, 16'd56727, 16'd61193, 16'd6197, 16'd55502, 16'd59258}; // indx = 3352
    #10;
    addra = 32'd107296;
    dina = {96'd0, 16'd65411, 16'd37890, 16'd30656, 16'd24963, 16'd19508, 16'd18231, 16'd56549, 16'd21588, 16'd15559, 16'd29627}; // indx = 3353
    #10;
    addra = 32'd107328;
    dina = {96'd0, 16'd10149, 16'd62139, 16'd41307, 16'd39401, 16'd65093, 16'd19889, 16'd6197, 16'd30774, 16'd2258, 16'd26655}; // indx = 3354
    #10;
    addra = 32'd107360;
    dina = {96'd0, 16'd6078, 16'd37804, 16'd5631, 16'd39457, 16'd47954, 16'd17484, 16'd30602, 16'd24503, 16'd33492, 16'd64973}; // indx = 3355
    #10;
    addra = 32'd107392;
    dina = {96'd0, 16'd48010, 16'd50561, 16'd64646, 16'd41070, 16'd4366, 16'd25107, 16'd52280, 16'd46855, 16'd26388, 16'd14317}; // indx = 3356
    #10;
    addra = 32'd107424;
    dina = {96'd0, 16'd44888, 16'd59899, 16'd21554, 16'd56010, 16'd39484, 16'd2461, 16'd11743, 16'd52236, 16'd41184, 16'd29931}; // indx = 3357
    #10;
    addra = 32'd107456;
    dina = {96'd0, 16'd21024, 16'd28509, 16'd38012, 16'd52868, 16'd55891, 16'd19944, 16'd29922, 16'd45284, 16'd17210, 16'd40312}; // indx = 3358
    #10;
    addra = 32'd107488;
    dina = {96'd0, 16'd11743, 16'd26625, 16'd64450, 16'd25220, 16'd51835, 16'd20645, 16'd16036, 16'd22618, 16'd50097, 16'd18005}; // indx = 3359
    #10;
    addra = 32'd107520;
    dina = {96'd0, 16'd62073, 16'd32818, 16'd39822, 16'd46144, 16'd30793, 16'd9661, 16'd26547, 16'd40718, 16'd17210, 16'd31495}; // indx = 3360
    #10;
    addra = 32'd107552;
    dina = {96'd0, 16'd10528, 16'd32343, 16'd46856, 16'd14309, 16'd58242, 16'd46102, 16'd36457, 16'd7331, 16'd5532, 16'd17201}; // indx = 3361
    #10;
    addra = 32'd107584;
    dina = {96'd0, 16'd53574, 16'd37105, 16'd13727, 16'd9879, 16'd18711, 16'd64711, 16'd31566, 16'd42801, 16'd56141, 16'd15319}; // indx = 3362
    #10;
    addra = 32'd107616;
    dina = {96'd0, 16'd47162, 16'd23826, 16'd21192, 16'd42074, 16'd24290, 16'd36689, 16'd15655, 16'd44780, 16'd46629, 16'd56968}; // indx = 3363
    #10;
    addra = 32'd107648;
    dina = {96'd0, 16'd48024, 16'd5531, 16'd837, 16'd11283, 16'd20998, 16'd12068, 16'd44659, 16'd33878, 16'd42365, 16'd27322}; // indx = 3364
    #10;
    addra = 32'd107680;
    dina = {96'd0, 16'd60123, 16'd38673, 16'd41304, 16'd55104, 16'd46692, 16'd53223, 16'd25432, 16'd46804, 16'd28493, 16'd36546}; // indx = 3365
    #10;
    addra = 32'd107712;
    dina = {96'd0, 16'd37971, 16'd54002, 16'd39309, 16'd23772, 16'd14995, 16'd60178, 16'd36928, 16'd46049, 16'd23819, 16'd40442}; // indx = 3366
    #10;
    addra = 32'd107744;
    dina = {96'd0, 16'd22613, 16'd42325, 16'd13056, 16'd47611, 16'd63015, 16'd18010, 16'd9708, 16'd27916, 16'd19484, 16'd12845}; // indx = 3367
    #10;
    addra = 32'd107776;
    dina = {96'd0, 16'd42098, 16'd32572, 16'd34666, 16'd48538, 16'd29744, 16'd7455, 16'd24964, 16'd42483, 16'd54985, 16'd58728}; // indx = 3368
    #10;
    addra = 32'd107808;
    dina = {96'd0, 16'd12824, 16'd15521, 16'd21513, 16'd32070, 16'd49010, 16'd21366, 16'd35784, 16'd13101, 16'd21896, 16'd28349}; // indx = 3369
    #10;
    addra = 32'd107840;
    dina = {96'd0, 16'd18763, 16'd7753, 16'd58510, 16'd25617, 16'd4574, 16'd56506, 16'd7833, 16'd23284, 16'd36738, 16'd22753}; // indx = 3370
    #10;
    addra = 32'd107872;
    dina = {96'd0, 16'd808, 16'd32615, 16'd57993, 16'd25982, 16'd39197, 16'd53693, 16'd8247, 16'd895, 16'd44633, 16'd39910}; // indx = 3371
    #10;
    addra = 32'd107904;
    dina = {96'd0, 16'd62658, 16'd44935, 16'd43829, 16'd23253, 16'd30562, 16'd65043, 16'd59698, 16'd31550, 16'd10739, 16'd20212}; // indx = 3372
    #10;
    addra = 32'd107936;
    dina = {96'd0, 16'd46244, 16'd31920, 16'd11152, 16'd10603, 16'd61165, 16'd33539, 16'd42706, 16'd381, 16'd60621, 16'd44280}; // indx = 3373
    #10;
    addra = 32'd107968;
    dina = {96'd0, 16'd64200, 16'd43898, 16'd59243, 16'd38354, 16'd42678, 16'd25204, 16'd79, 16'd167, 16'd2151, 16'd2816}; // indx = 3374
    #10;
    addra = 32'd108000;
    dina = {96'd0, 16'd43604, 16'd20671, 16'd32475, 16'd36681, 16'd49004, 16'd36689, 16'd38288, 16'd15575, 16'd65142, 16'd61065}; // indx = 3375
    #10;
    addra = 32'd108032;
    dina = {96'd0, 16'd43948, 16'd4192, 16'd53425, 16'd50661, 16'd13396, 16'd22017, 16'd54088, 16'd60340, 16'd49384, 16'd60070}; // indx = 3376
    #10;
    addra = 32'd108064;
    dina = {96'd0, 16'd38829, 16'd15667, 16'd33792, 16'd8856, 16'd32984, 16'd26507, 16'd22744, 16'd33922, 16'd62488, 16'd62018}; // indx = 3377
    #10;
    addra = 32'd108096;
    dina = {96'd0, 16'd27192, 16'd45167, 16'd54592, 16'd45555, 16'd56723, 16'd40434, 16'd5238, 16'd40212, 16'd16590, 16'd54942}; // indx = 3378
    #10;
    addra = 32'd108128;
    dina = {96'd0, 16'd22778, 16'd5191, 16'd43644, 16'd18759, 16'd35843, 16'd43394, 16'd60701, 16'd26256, 16'd12197, 16'd63790}; // indx = 3379
    #10;
    addra = 32'd108160;
    dina = {96'd0, 16'd48722, 16'd46046, 16'd33918, 16'd53610, 16'd3320, 16'd7331, 16'd20760, 16'd56314, 16'd43487, 16'd58588}; // indx = 3380
    #10;
    addra = 32'd108192;
    dina = {96'd0, 16'd40344, 16'd42667, 16'd44899, 16'd28386, 16'd11106, 16'd26046, 16'd42286, 16'd11288, 16'd18859, 16'd46913}; // indx = 3381
    #10;
    addra = 32'd108224;
    dina = {96'd0, 16'd16167, 16'd41554, 16'd31116, 16'd61049, 16'd50153, 16'd1464, 16'd2901, 16'd40831, 16'd48506, 16'd22695}; // indx = 3382
    #10;
    addra = 32'd108256;
    dina = {96'd0, 16'd57733, 16'd56311, 16'd29221, 16'd42586, 16'd39078, 16'd27156, 16'd46117, 16'd37263, 16'd16629, 16'd52332}; // indx = 3383
    #10;
    addra = 32'd108288;
    dina = {96'd0, 16'd48803, 16'd35345, 16'd36301, 16'd22025, 16'd48049, 16'd31571, 16'd63205, 16'd65334, 16'd59813, 16'd60237}; // indx = 3384
    #10;
    addra = 32'd108320;
    dina = {96'd0, 16'd10020, 16'd46810, 16'd48048, 16'd56756, 16'd24342, 16'd38917, 16'd18696, 16'd44916, 16'd9363, 16'd349}; // indx = 3385
    #10;
    addra = 32'd108352;
    dina = {96'd0, 16'd6974, 16'd9421, 16'd27341, 16'd64791, 16'd3922, 16'd45479, 16'd9389, 16'd15410, 16'd23298, 16'd6004}; // indx = 3386
    #10;
    addra = 32'd108384;
    dina = {96'd0, 16'd37421, 16'd46256, 16'd33938, 16'd5990, 16'd45279, 16'd55747, 16'd41477, 16'd62868, 16'd21731, 16'd33286}; // indx = 3387
    #10;
    addra = 32'd108416;
    dina = {96'd0, 16'd4734, 16'd23761, 16'd52384, 16'd48127, 16'd13535, 16'd1357, 16'd32985, 16'd12366, 16'd9508, 16'd19095}; // indx = 3388
    #10;
    addra = 32'd108448;
    dina = {96'd0, 16'd59289, 16'd62499, 16'd28364, 16'd30196, 16'd23840, 16'd16269, 16'd5404, 16'd45984, 16'd9558, 16'd34488}; // indx = 3389
    #10;
    addra = 32'd108480;
    dina = {96'd0, 16'd27388, 16'd36522, 16'd56447, 16'd21029, 16'd10935, 16'd3488, 16'd11356, 16'd59999, 16'd10324, 16'd58362}; // indx = 3390
    #10;
    addra = 32'd108512;
    dina = {96'd0, 16'd28024, 16'd46907, 16'd21027, 16'd10507, 16'd41775, 16'd32563, 16'd48629, 16'd63272, 16'd37971, 16'd30571}; // indx = 3391
    #10;
    addra = 32'd108544;
    dina = {96'd0, 16'd45778, 16'd36063, 16'd21888, 16'd52324, 16'd7449, 16'd28906, 16'd46188, 16'd37707, 16'd47405, 16'd19065}; // indx = 3392
    #10;
    addra = 32'd108576;
    dina = {96'd0, 16'd47187, 16'd44483, 16'd21228, 16'd56725, 16'd62291, 16'd17457, 16'd11715, 16'd59218, 16'd20977, 16'd23602}; // indx = 3393
    #10;
    addra = 32'd108608;
    dina = {96'd0, 16'd29562, 16'd5655, 16'd39806, 16'd20628, 16'd39921, 16'd29382, 16'd28198, 16'd24722, 16'd9144, 16'd22256}; // indx = 3394
    #10;
    addra = 32'd108640;
    dina = {96'd0, 16'd40127, 16'd17386, 16'd17337, 16'd52987, 16'd48712, 16'd45483, 16'd65167, 16'd32207, 16'd50907, 16'd1286}; // indx = 3395
    #10;
    addra = 32'd108672;
    dina = {96'd0, 16'd55225, 16'd41119, 16'd63050, 16'd15443, 16'd60611, 16'd3501, 16'd52167, 16'd62898, 16'd64156, 16'd56702}; // indx = 3396
    #10;
    addra = 32'd108704;
    dina = {96'd0, 16'd45564, 16'd17919, 16'd47435, 16'd13090, 16'd53056, 16'd57017, 16'd18187, 16'd26633, 16'd33605, 16'd11179}; // indx = 3397
    #10;
    addra = 32'd108736;
    dina = {96'd0, 16'd50015, 16'd32680, 16'd28956, 16'd17978, 16'd45378, 16'd13977, 16'd9336, 16'd15181, 16'd2614, 16'd63664}; // indx = 3398
    #10;
    addra = 32'd108768;
    dina = {96'd0, 16'd62676, 16'd19156, 16'd42657, 16'd58344, 16'd51598, 16'd14047, 16'd63571, 16'd49250, 16'd2997, 16'd63973}; // indx = 3399
    #10;
    addra = 32'd108800;
    dina = {96'd0, 16'd26832, 16'd13612, 16'd59162, 16'd26907, 16'd43415, 16'd19986, 16'd48688, 16'd23708, 16'd2315, 16'd11056}; // indx = 3400
    #10;
    addra = 32'd108832;
    dina = {96'd0, 16'd28749, 16'd5631, 16'd1666, 16'd62355, 16'd37087, 16'd12795, 16'd26000, 16'd47657, 16'd21064, 16'd4688}; // indx = 3401
    #10;
    addra = 32'd108864;
    dina = {96'd0, 16'd29595, 16'd46732, 16'd22565, 16'd21768, 16'd52798, 16'd43326, 16'd1576, 16'd14011, 16'd30416, 16'd27643}; // indx = 3402
    #10;
    addra = 32'd108896;
    dina = {96'd0, 16'd58869, 16'd48956, 16'd2740, 16'd21057, 16'd4451, 16'd34932, 16'd53760, 16'd10220, 16'd23664, 16'd15017}; // indx = 3403
    #10;
    addra = 32'd108928;
    dina = {96'd0, 16'd35913, 16'd46667, 16'd2282, 16'd2840, 16'd20538, 16'd20422, 16'd61293, 16'd45668, 16'd51728, 16'd6228}; // indx = 3404
    #10;
    addra = 32'd108960;
    dina = {96'd0, 16'd56199, 16'd33598, 16'd39995, 16'd13089, 16'd1045, 16'd12430, 16'd39858, 16'd16895, 16'd51530, 16'd41087}; // indx = 3405
    #10;
    addra = 32'd108992;
    dina = {96'd0, 16'd12338, 16'd14055, 16'd1147, 16'd25033, 16'd31916, 16'd26259, 16'd3566, 16'd3433, 16'd20793, 16'd35723}; // indx = 3406
    #10;
    addra = 32'd109024;
    dina = {96'd0, 16'd4435, 16'd36182, 16'd39741, 16'd2203, 16'd34488, 16'd46926, 16'd42388, 16'd2972, 16'd47676, 16'd10954}; // indx = 3407
    #10;
    addra = 32'd109056;
    dina = {96'd0, 16'd38946, 16'd42289, 16'd44076, 16'd38491, 16'd35993, 16'd23235, 16'd6672, 16'd60671, 16'd45491, 16'd24895}; // indx = 3408
    #10;
    addra = 32'd109088;
    dina = {96'd0, 16'd50877, 16'd56911, 16'd14378, 16'd2636, 16'd53637, 16'd40190, 16'd58898, 16'd13138, 16'd4211, 16'd59465}; // indx = 3409
    #10;
    addra = 32'd109120;
    dina = {96'd0, 16'd33213, 16'd59371, 16'd11266, 16'd27210, 16'd63145, 16'd24063, 16'd64616, 16'd5885, 16'd48629, 16'd40868}; // indx = 3410
    #10;
    addra = 32'd109152;
    dina = {96'd0, 16'd51041, 16'd64453, 16'd12465, 16'd37908, 16'd22031, 16'd1620, 16'd29848, 16'd46345, 16'd63004, 16'd29732}; // indx = 3411
    #10;
    addra = 32'd109184;
    dina = {96'd0, 16'd46909, 16'd3648, 16'd1869, 16'd463, 16'd59451, 16'd2685, 16'd2761, 16'd10326, 16'd29536, 16'd62728}; // indx = 3412
    #10;
    addra = 32'd109216;
    dina = {96'd0, 16'd9014, 16'd47287, 16'd34615, 16'd59236, 16'd39982, 16'd20599, 16'd27132, 16'd9079, 16'd46705, 16'd64379}; // indx = 3413
    #10;
    addra = 32'd109248;
    dina = {96'd0, 16'd45800, 16'd32671, 16'd20037, 16'd46684, 16'd62353, 16'd19460, 16'd62293, 16'd64383, 16'd24640, 16'd199}; // indx = 3414
    #10;
    addra = 32'd109280;
    dina = {96'd0, 16'd55923, 16'd54078, 16'd33257, 16'd55010, 16'd3031, 16'd49656, 16'd59761, 16'd51848, 16'd52086, 16'd25489}; // indx = 3415
    #10;
    addra = 32'd109312;
    dina = {96'd0, 16'd28320, 16'd21326, 16'd54194, 16'd15668, 16'd53301, 16'd9645, 16'd57383, 16'd34212, 16'd50321, 16'd33515}; // indx = 3416
    #10;
    addra = 32'd109344;
    dina = {96'd0, 16'd40872, 16'd41852, 16'd22886, 16'd54243, 16'd28590, 16'd37838, 16'd15733, 16'd58892, 16'd54412, 16'd55695}; // indx = 3417
    #10;
    addra = 32'd109376;
    dina = {96'd0, 16'd43977, 16'd48916, 16'd36312, 16'd5936, 16'd54122, 16'd58932, 16'd39816, 16'd36132, 16'd36791, 16'd47293}; // indx = 3418
    #10;
    addra = 32'd109408;
    dina = {96'd0, 16'd13800, 16'd37856, 16'd63412, 16'd36932, 16'd59662, 16'd27308, 16'd62959, 16'd36988, 16'd42567, 16'd49869}; // indx = 3419
    #10;
    addra = 32'd109440;
    dina = {96'd0, 16'd2896, 16'd51230, 16'd36054, 16'd30454, 16'd21378, 16'd58928, 16'd57438, 16'd64474, 16'd17859, 16'd21665}; // indx = 3420
    #10;
    addra = 32'd109472;
    dina = {96'd0, 16'd56854, 16'd1450, 16'd635, 16'd59609, 16'd63205, 16'd44427, 16'd15563, 16'd53310, 16'd21263, 16'd10583}; // indx = 3421
    #10;
    addra = 32'd109504;
    dina = {96'd0, 16'd52743, 16'd30947, 16'd19487, 16'd22317, 16'd12134, 16'd31280, 16'd61334, 16'd59416, 16'd26251, 16'd39773}; // indx = 3422
    #10;
    addra = 32'd109536;
    dina = {96'd0, 16'd30176, 16'd63947, 16'd28071, 16'd6375, 16'd24434, 16'd15494, 16'd9925, 16'd21695, 16'd15744, 16'd6338}; // indx = 3423
    #10;
    addra = 32'd109568;
    dina = {96'd0, 16'd24335, 16'd2616, 16'd4414, 16'd15756, 16'd55297, 16'd17700, 16'd46529, 16'd58667, 16'd10163, 16'd16736}; // indx = 3424
    #10;
    addra = 32'd109600;
    dina = {96'd0, 16'd48928, 16'd28246, 16'd38194, 16'd63335, 16'd41327, 16'd177, 16'd23671, 16'd45189, 16'd61882, 16'd14237}; // indx = 3425
    #10;
    addra = 32'd109632;
    dina = {96'd0, 16'd39383, 16'd55185, 16'd30691, 16'd39720, 16'd20877, 16'd59062, 16'd46377, 16'd52809, 16'd285, 16'd45671}; // indx = 3426
    #10;
    addra = 32'd109664;
    dina = {96'd0, 16'd46728, 16'd26579, 16'd41301, 16'd36827, 16'd64173, 16'd17707, 16'd16234, 16'd64855, 16'd11759, 16'd5858}; // indx = 3427
    #10;
    addra = 32'd109696;
    dina = {96'd0, 16'd40325, 16'd28769, 16'd49496, 16'd14487, 16'd36856, 16'd62388, 16'd55253, 16'd63618, 16'd16589, 16'd51320}; // indx = 3428
    #10;
    addra = 32'd109728;
    dina = {96'd0, 16'd63267, 16'd14462, 16'd2230, 16'd42095, 16'd57700, 16'd3698, 16'd30101, 16'd27303, 16'd30336, 16'd59374}; // indx = 3429
    #10;
    addra = 32'd109760;
    dina = {96'd0, 16'd61618, 16'd42297, 16'd17962, 16'd33421, 16'd55650, 16'd4244, 16'd18628, 16'd46527, 16'd35972, 16'd19787}; // indx = 3430
    #10;
    addra = 32'd109792;
    dina = {96'd0, 16'd43679, 16'd19109, 16'd56606, 16'd40712, 16'd29342, 16'd2172, 16'd58436, 16'd45253, 16'd16239, 16'd61519}; // indx = 3431
    #10;
    addra = 32'd109824;
    dina = {96'd0, 16'd38009, 16'd39562, 16'd2003, 16'd31172, 16'd30061, 16'd18403, 16'd3671, 16'd48128, 16'd51448, 16'd48815}; // indx = 3432
    #10;
    addra = 32'd109856;
    dina = {96'd0, 16'd11893, 16'd21681, 16'd47406, 16'd64476, 16'd26946, 16'd9217, 16'd50100, 16'd360, 16'd44905, 16'd64530}; // indx = 3433
    #10;
    addra = 32'd109888;
    dina = {96'd0, 16'd56171, 16'd48283, 16'd14369, 16'd57319, 16'd48708, 16'd47526, 16'd61139, 16'd30535, 16'd34254, 16'd3252}; // indx = 3434
    #10;
    addra = 32'd109920;
    dina = {96'd0, 16'd24876, 16'd58530, 16'd3641, 16'd13582, 16'd39280, 16'd64384, 16'd17669, 16'd38968, 16'd24477, 16'd25392}; // indx = 3435
    #10;
    addra = 32'd109952;
    dina = {96'd0, 16'd30038, 16'd40196, 16'd52691, 16'd24338, 16'd40027, 16'd65368, 16'd14001, 16'd19097, 16'd33558, 16'd51686}; // indx = 3436
    #10;
    addra = 32'd109984;
    dina = {96'd0, 16'd39070, 16'd55595, 16'd65154, 16'd41802, 16'd56538, 16'd59632, 16'd62056, 16'd63269, 16'd53870, 16'd62429}; // indx = 3437
    #10;
    addra = 32'd110016;
    dina = {96'd0, 16'd56185, 16'd11489, 16'd43519, 16'd44840, 16'd7352, 16'd8776, 16'd31399, 16'd60984, 16'd28238, 16'd34281}; // indx = 3438
    #10;
    addra = 32'd110048;
    dina = {96'd0, 16'd3440, 16'd35767, 16'd22325, 16'd34844, 16'd20814, 16'd5986, 16'd59869, 16'd61741, 16'd64842, 16'd31920}; // indx = 3439
    #10;
    addra = 32'd110080;
    dina = {96'd0, 16'd25838, 16'd30878, 16'd7669, 16'd41415, 16'd26482, 16'd48861, 16'd31072, 16'd29276, 16'd24305, 16'd1950}; // indx = 3440
    #10;
    addra = 32'd110112;
    dina = {96'd0, 16'd58589, 16'd44568, 16'd10092, 16'd34135, 16'd60687, 16'd29951, 16'd25903, 16'd33547, 16'd15426, 16'd32044}; // indx = 3441
    #10;
    addra = 32'd110144;
    dina = {96'd0, 16'd59570, 16'd39528, 16'd48395, 16'd19853, 16'd15560, 16'd34035, 16'd10428, 16'd24076, 16'd52880, 16'd36254}; // indx = 3442
    #10;
    addra = 32'd110176;
    dina = {96'd0, 16'd34343, 16'd26315, 16'd65413, 16'd14659, 16'd43303, 16'd40342, 16'd18231, 16'd9140, 16'd27664, 16'd5549}; // indx = 3443
    #10;
    addra = 32'd110208;
    dina = {96'd0, 16'd23604, 16'd22861, 16'd17555, 16'd41519, 16'd35259, 16'd5653, 16'd8468, 16'd534, 16'd43150, 16'd45660}; // indx = 3444
    #10;
    addra = 32'd110240;
    dina = {96'd0, 16'd56803, 16'd7571, 16'd38947, 16'd56593, 16'd45574, 16'd30695, 16'd15409, 16'd61218, 16'd8848, 16'd64217}; // indx = 3445
    #10;
    addra = 32'd110272;
    dina = {96'd0, 16'd47910, 16'd21958, 16'd57808, 16'd4288, 16'd54348, 16'd17669, 16'd28667, 16'd48155, 16'd40189, 16'd45577}; // indx = 3446
    #10;
    addra = 32'd110304;
    dina = {96'd0, 16'd1664, 16'd21386, 16'd2453, 16'd35347, 16'd58999, 16'd60418, 16'd25068, 16'd7541, 16'd40326, 16'd41417}; // indx = 3447
    #10;
    addra = 32'd110336;
    dina = {96'd0, 16'd9922, 16'd50944, 16'd14625, 16'd57013, 16'd19994, 16'd53266, 16'd23785, 16'd59222, 16'd45952, 16'd56980}; // indx = 3448
    #10;
    addra = 32'd110368;
    dina = {96'd0, 16'd6281, 16'd35210, 16'd42086, 16'd58431, 16'd6825, 16'd60182, 16'd63887, 16'd37312, 16'd3767, 16'd58087}; // indx = 3449
    #10;
    addra = 32'd110400;
    dina = {96'd0, 16'd30027, 16'd37377, 16'd41647, 16'd32043, 16'd30520, 16'd6329, 16'd47794, 16'd33991, 16'd54720, 16'd1182}; // indx = 3450
    #10;
    addra = 32'd110432;
    dina = {96'd0, 16'd12177, 16'd15413, 16'd5901, 16'd56808, 16'd56559, 16'd62883, 16'd18606, 16'd63982, 16'd11553, 16'd1716}; // indx = 3451
    #10;
    addra = 32'd110464;
    dina = {96'd0, 16'd4920, 16'd46396, 16'd23300, 16'd33882, 16'd48589, 16'd35648, 16'd17554, 16'd51573, 16'd11847, 16'd27591}; // indx = 3452
    #10;
    addra = 32'd110496;
    dina = {96'd0, 16'd14606, 16'd8623, 16'd33659, 16'd54509, 16'd59576, 16'd38067, 16'd43294, 16'd408, 16'd58289, 16'd26325}; // indx = 3453
    #10;
    addra = 32'd110528;
    dina = {96'd0, 16'd60138, 16'd5390, 16'd31324, 16'd44874, 16'd24924, 16'd65026, 16'd21198, 16'd12351, 16'd40230, 16'd8144}; // indx = 3454
    #10;
    addra = 32'd110560;
    dina = {96'd0, 16'd27936, 16'd4570, 16'd30459, 16'd62665, 16'd15166, 16'd54449, 16'd3247, 16'd35014, 16'd14474, 16'd34889}; // indx = 3455
    #10;
    addra = 32'd110592;
    dina = {96'd0, 16'd47256, 16'd62265, 16'd6114, 16'd16863, 16'd26139, 16'd54463, 16'd54882, 16'd2231, 16'd40852, 16'd43045}; // indx = 3456
    #10;
    addra = 32'd110624;
    dina = {96'd0, 16'd33558, 16'd52950, 16'd17322, 16'd23300, 16'd48884, 16'd47093, 16'd33377, 16'd88, 16'd47408, 16'd39465}; // indx = 3457
    #10;
    addra = 32'd110656;
    dina = {96'd0, 16'd60959, 16'd4626, 16'd40731, 16'd60671, 16'd50960, 16'd58312, 16'd53421, 16'd23596, 16'd63975, 16'd15480}; // indx = 3458
    #10;
    addra = 32'd110688;
    dina = {96'd0, 16'd65242, 16'd46784, 16'd31989, 16'd29684, 16'd5695, 16'd33012, 16'd3155, 16'd48663, 16'd25227, 16'd52742}; // indx = 3459
    #10;
    addra = 32'd110720;
    dina = {96'd0, 16'd62641, 16'd51565, 16'd29493, 16'd55998, 16'd30771, 16'd65246, 16'd22212, 16'd44827, 16'd13443, 16'd24484}; // indx = 3460
    #10;
    addra = 32'd110752;
    dina = {96'd0, 16'd16667, 16'd43342, 16'd31405, 16'd19488, 16'd3852, 16'd49278, 16'd42977, 16'd15948, 16'd34554, 16'd21214}; // indx = 3461
    #10;
    addra = 32'd110784;
    dina = {96'd0, 16'd50938, 16'd49036, 16'd49959, 16'd28241, 16'd19209, 16'd28447, 16'd33473, 16'd30045, 16'd6806, 16'd25633}; // indx = 3462
    #10;
    addra = 32'd110816;
    dina = {96'd0, 16'd29870, 16'd6848, 16'd19526, 16'd20640, 16'd43364, 16'd15892, 16'd55222, 16'd966, 16'd40210, 16'd48270}; // indx = 3463
    #10;
    addra = 32'd110848;
    dina = {96'd0, 16'd57202, 16'd55427, 16'd2406, 16'd46696, 16'd32144, 16'd59428, 16'd50803, 16'd55113, 16'd2382, 16'd33816}; // indx = 3464
    #10;
    addra = 32'd110880;
    dina = {96'd0, 16'd6966, 16'd3365, 16'd63033, 16'd11386, 16'd41596, 16'd9966, 16'd46651, 16'd38782, 16'd20686, 16'd60750}; // indx = 3465
    #10;
    addra = 32'd110912;
    dina = {96'd0, 16'd15491, 16'd29679, 16'd28716, 16'd14065, 16'd6264, 16'd21499, 16'd40150, 16'd46417, 16'd56451, 16'd32647}; // indx = 3466
    #10;
    addra = 32'd110944;
    dina = {96'd0, 16'd39575, 16'd19051, 16'd26207, 16'd45590, 16'd56779, 16'd12984, 16'd8084, 16'd1172, 16'd23855, 16'd50631}; // indx = 3467
    #10;
    addra = 32'd110976;
    dina = {96'd0, 16'd43497, 16'd24171, 16'd54586, 16'd52961, 16'd26400, 16'd28264, 16'd19359, 16'd10337, 16'd34907, 16'd28149}; // indx = 3468
    #10;
    addra = 32'd111008;
    dina = {96'd0, 16'd13658, 16'd41765, 16'd13592, 16'd63950, 16'd47407, 16'd15959, 16'd38414, 16'd59460, 16'd25384, 16'd30352}; // indx = 3469
    #10;
    addra = 32'd111040;
    dina = {96'd0, 16'd60611, 16'd31876, 16'd20692, 16'd33940, 16'd27213, 16'd63230, 16'd19770, 16'd36189, 16'd13412, 16'd62194}; // indx = 3470
    #10;
    addra = 32'd111072;
    dina = {96'd0, 16'd62071, 16'd3319, 16'd39178, 16'd40601, 16'd21650, 16'd46372, 16'd14342, 16'd36152, 16'd7639, 16'd22197}; // indx = 3471
    #10;
    addra = 32'd111104;
    dina = {96'd0, 16'd59022, 16'd18219, 16'd22832, 16'd24239, 16'd20684, 16'd19686, 16'd1101, 16'd24938, 16'd64780, 16'd40259}; // indx = 3472
    #10;
    addra = 32'd111136;
    dina = {96'd0, 16'd51296, 16'd18501, 16'd60811, 16'd27938, 16'd9329, 16'd49081, 16'd6871, 16'd26315, 16'd40447, 16'd30240}; // indx = 3473
    #10;
    addra = 32'd111168;
    dina = {96'd0, 16'd55950, 16'd44665, 16'd26400, 16'd35494, 16'd60262, 16'd32613, 16'd11571, 16'd15543, 16'd45123, 16'd58203}; // indx = 3474
    #10;
    addra = 32'd111200;
    dina = {96'd0, 16'd19812, 16'd5295, 16'd8424, 16'd15406, 16'd32900, 16'd23566, 16'd29302, 16'd64251, 16'd27807, 16'd48002}; // indx = 3475
    #10;
    addra = 32'd111232;
    dina = {96'd0, 16'd38710, 16'd49349, 16'd57136, 16'd14562, 16'd51425, 16'd14332, 16'd16441, 16'd35357, 16'd48929, 16'd63523}; // indx = 3476
    #10;
    addra = 32'd111264;
    dina = {96'd0, 16'd59830, 16'd7528, 16'd4842, 16'd50427, 16'd40890, 16'd41213, 16'd19247, 16'd12709, 16'd9888, 16'd61217}; // indx = 3477
    #10;
    addra = 32'd111296;
    dina = {96'd0, 16'd1819, 16'd26995, 16'd43124, 16'd54270, 16'd11542, 16'd26963, 16'd54663, 16'd8127, 16'd58038, 16'd11540}; // indx = 3478
    #10;
    addra = 32'd111328;
    dina = {96'd0, 16'd22, 16'd19970, 16'd38921, 16'd6065, 16'd21554, 16'd6728, 16'd9451, 16'd21858, 16'd37256, 16'd26074}; // indx = 3479
    #10;
    addra = 32'd111360;
    dina = {96'd0, 16'd16054, 16'd40556, 16'd48689, 16'd6047, 16'd46971, 16'd5840, 16'd9126, 16'd31100, 16'd52519, 16'd2239}; // indx = 3480
    #10;
    addra = 32'd111392;
    dina = {96'd0, 16'd42412, 16'd31591, 16'd52193, 16'd27608, 16'd43539, 16'd41747, 16'd64967, 16'd65348, 16'd65388, 16'd29277}; // indx = 3481
    #10;
    addra = 32'd111424;
    dina = {96'd0, 16'd3733, 16'd51250, 16'd24629, 16'd24239, 16'd19476, 16'd46622, 16'd49391, 16'd18616, 16'd19659, 16'd3673}; // indx = 3482
    #10;
    addra = 32'd111456;
    dina = {96'd0, 16'd54435, 16'd31265, 16'd56197, 16'd32726, 16'd29467, 16'd10524, 16'd3999, 16'd2620, 16'd44880, 16'd63466}; // indx = 3483
    #10;
    addra = 32'd111488;
    dina = {96'd0, 16'd54383, 16'd54923, 16'd19951, 16'd24942, 16'd21133, 16'd49401, 16'd18897, 16'd56357, 16'd36281, 16'd37875}; // indx = 3484
    #10;
    addra = 32'd111520;
    dina = {96'd0, 16'd9766, 16'd3777, 16'd40951, 16'd7770, 16'd4681, 16'd20739, 16'd5108, 16'd63303, 16'd29710, 16'd43059}; // indx = 3485
    #10;
    addra = 32'd111552;
    dina = {96'd0, 16'd3046, 16'd27510, 16'd63231, 16'd35004, 16'd58024, 16'd50712, 16'd2442, 16'd36624, 16'd5784, 16'd18559}; // indx = 3486
    #10;
    addra = 32'd111584;
    dina = {96'd0, 16'd41501, 16'd63428, 16'd39712, 16'd43229, 16'd20336, 16'd21220, 16'd14447, 16'd39362, 16'd23824, 16'd62880}; // indx = 3487
    #10;
    addra = 32'd111616;
    dina = {96'd0, 16'd63786, 16'd60258, 16'd47114, 16'd31430, 16'd28271, 16'd46568, 16'd41071, 16'd36275, 16'd53121, 16'd46047}; // indx = 3488
    #10;
    addra = 32'd111648;
    dina = {96'd0, 16'd10999, 16'd24023, 16'd60944, 16'd52247, 16'd63935, 16'd5136, 16'd57122, 16'd12641, 16'd36444, 16'd39202}; // indx = 3489
    #10;
    addra = 32'd111680;
    dina = {96'd0, 16'd31228, 16'd26006, 16'd5213, 16'd57877, 16'd34924, 16'd39036, 16'd115, 16'd34446, 16'd27766, 16'd61386}; // indx = 3490
    #10;
    addra = 32'd111712;
    dina = {96'd0, 16'd52276, 16'd17465, 16'd819, 16'd30520, 16'd40923, 16'd12142, 16'd24090, 16'd9585, 16'd44002, 16'd39430}; // indx = 3491
    #10;
    addra = 32'd111744;
    dina = {96'd0, 16'd28983, 16'd11632, 16'd53316, 16'd60069, 16'd48624, 16'd1148, 16'd9936, 16'd43274, 16'd20771, 16'd7524}; // indx = 3492
    #10;
    addra = 32'd111776;
    dina = {96'd0, 16'd44698, 16'd46417, 16'd19392, 16'd15539, 16'd6777, 16'd20235, 16'd29326, 16'd22201, 16'd14677, 16'd30814}; // indx = 3493
    #10;
    addra = 32'd111808;
    dina = {96'd0, 16'd62620, 16'd1066, 16'd16849, 16'd4910, 16'd13957, 16'd38585, 16'd13466, 16'd51562, 16'd23225, 16'd17704}; // indx = 3494
    #10;
    addra = 32'd111840;
    dina = {96'd0, 16'd44667, 16'd36326, 16'd7588, 16'd13406, 16'd50606, 16'd45871, 16'd23263, 16'd23933, 16'd16226, 16'd23287}; // indx = 3495
    #10;
    addra = 32'd111872;
    dina = {96'd0, 16'd30421, 16'd32576, 16'd14545, 16'd30443, 16'd36194, 16'd56408, 16'd22763, 16'd17050, 16'd49925, 16'd2358}; // indx = 3496
    #10;
    addra = 32'd111904;
    dina = {96'd0, 16'd38143, 16'd45138, 16'd2493, 16'd4183, 16'd46813, 16'd25794, 16'd26082, 16'd59558, 16'd34316, 16'd18180}; // indx = 3497
    #10;
    addra = 32'd111936;
    dina = {96'd0, 16'd24661, 16'd26948, 16'd11012, 16'd11828, 16'd1716, 16'd39637, 16'd21126, 16'd60245, 16'd43243, 16'd58364}; // indx = 3498
    #10;
    addra = 32'd111968;
    dina = {96'd0, 16'd58161, 16'd24558, 16'd25676, 16'd6379, 16'd49512, 16'd20499, 16'd37867, 16'd26767, 16'd36374, 16'd58417}; // indx = 3499
    #10;
    addra = 32'd112000;
    dina = {96'd0, 16'd61534, 16'd3392, 16'd36459, 16'd34559, 16'd40167, 16'd40568, 16'd30351, 16'd26517, 16'd62117, 16'd43034}; // indx = 3500
    #10;
    addra = 32'd112032;
    dina = {96'd0, 16'd14906, 16'd50276, 16'd3224, 16'd21556, 16'd20404, 16'd34897, 16'd47237, 16'd14842, 16'd56780, 16'd28710}; // indx = 3501
    #10;
    addra = 32'd112064;
    dina = {96'd0, 16'd14169, 16'd20416, 16'd2334, 16'd20510, 16'd57966, 16'd44868, 16'd9472, 16'd27389, 16'd1964, 16'd65452}; // indx = 3502
    #10;
    addra = 32'd112096;
    dina = {96'd0, 16'd3177, 16'd49567, 16'd47457, 16'd19044, 16'd41926, 16'd8589, 16'd29802, 16'd22822, 16'd29849, 16'd12959}; // indx = 3503
    #10;
    addra = 32'd112128;
    dina = {96'd0, 16'd21071, 16'd57491, 16'd11159, 16'd34153, 16'd46512, 16'd11828, 16'd32001, 16'd671, 16'd13116, 16'd19532}; // indx = 3504
    #10;
    addra = 32'd112160;
    dina = {96'd0, 16'd52732, 16'd50349, 16'd25038, 16'd41977, 16'd41704, 16'd55987, 16'd54311, 16'd24922, 16'd36054, 16'd43431}; // indx = 3505
    #10;
    addra = 32'd112192;
    dina = {96'd0, 16'd18177, 16'd46364, 16'd62921, 16'd49422, 16'd15298, 16'd14758, 16'd33181, 16'd43565, 16'd60429, 16'd19309}; // indx = 3506
    #10;
    addra = 32'd112224;
    dina = {96'd0, 16'd42496, 16'd49061, 16'd29605, 16'd21168, 16'd36306, 16'd2761, 16'd36599, 16'd57688, 16'd56904, 16'd27672}; // indx = 3507
    #10;
    addra = 32'd112256;
    dina = {96'd0, 16'd50259, 16'd60672, 16'd56537, 16'd33921, 16'd45101, 16'd42564, 16'd790, 16'd61194, 16'd14787, 16'd22994}; // indx = 3508
    #10;
    addra = 32'd112288;
    dina = {96'd0, 16'd19869, 16'd14155, 16'd13441, 16'd8515, 16'd31083, 16'd64200, 16'd46922, 16'd23200, 16'd29076, 16'd12296}; // indx = 3509
    #10;
    addra = 32'd112320;
    dina = {96'd0, 16'd39962, 16'd6152, 16'd34937, 16'd48752, 16'd11238, 16'd86, 16'd34195, 16'd50079, 16'd34498, 16'd2364}; // indx = 3510
    #10;
    addra = 32'd112352;
    dina = {96'd0, 16'd12529, 16'd25635, 16'd45632, 16'd63335, 16'd4673, 16'd36495, 16'd21750, 16'd11638, 16'd4464, 16'd34698}; // indx = 3511
    #10;
    addra = 32'd112384;
    dina = {96'd0, 16'd3222, 16'd41199, 16'd29760, 16'd9749, 16'd17166, 16'd5723, 16'd17133, 16'd19315, 16'd34737, 16'd41315}; // indx = 3512
    #10;
    addra = 32'd112416;
    dina = {96'd0, 16'd3045, 16'd29094, 16'd6382, 16'd18829, 16'd41959, 16'd54528, 16'd58340, 16'd22259, 16'd36527, 16'd44380}; // indx = 3513
    #10;
    addra = 32'd112448;
    dina = {96'd0, 16'd41309, 16'd20147, 16'd20642, 16'd50890, 16'd15975, 16'd53846, 16'd40866, 16'd60303, 16'd46597, 16'd61538}; // indx = 3514
    #10;
    addra = 32'd112480;
    dina = {96'd0, 16'd4158, 16'd41726, 16'd23415, 16'd27565, 16'd4953, 16'd57414, 16'd62253, 16'd31691, 16'd36128, 16'd26195}; // indx = 3515
    #10;
    addra = 32'd112512;
    dina = {96'd0, 16'd22493, 16'd36575, 16'd63332, 16'd36118, 16'd20076, 16'd16049, 16'd20969, 16'd21659, 16'd27720, 16'd60333}; // indx = 3516
    #10;
    addra = 32'd112544;
    dina = {96'd0, 16'd2894, 16'd46259, 16'd51131, 16'd50117, 16'd2712, 16'd44815, 16'd17471, 16'd445, 16'd50698, 16'd46692}; // indx = 3517
    #10;
    addra = 32'd112576;
    dina = {96'd0, 16'd16178, 16'd30245, 16'd51595, 16'd22937, 16'd22937, 16'd54273, 16'd28849, 16'd34963, 16'd54048, 16'd20385}; // indx = 3518
    #10;
    addra = 32'd112608;
    dina = {96'd0, 16'd63424, 16'd9341, 16'd29199, 16'd37400, 16'd50480, 16'd64580, 16'd2395, 16'd26439, 16'd56887, 16'd11099}; // indx = 3519
    #10;
    addra = 32'd112640;
    dina = {96'd0, 16'd45364, 16'd16868, 16'd35877, 16'd16068, 16'd37983, 16'd24131, 16'd266, 16'd12743, 16'd21717, 16'd25745}; // indx = 3520
    #10;
    addra = 32'd112672;
    dina = {96'd0, 16'd53663, 16'd42917, 16'd63754, 16'd63266, 16'd8114, 16'd37663, 16'd50803, 16'd4877, 16'd38786, 16'd11804}; // indx = 3521
    #10;
    addra = 32'd112704;
    dina = {96'd0, 16'd60218, 16'd55992, 16'd45429, 16'd12803, 16'd22042, 16'd59631, 16'd49639, 16'd53484, 16'd59526, 16'd63631}; // indx = 3522
    #10;
    addra = 32'd112736;
    dina = {96'd0, 16'd29721, 16'd29862, 16'd16478, 16'd19167, 16'd2266, 16'd23115, 16'd2579, 16'd35729, 16'd27162, 16'd25768}; // indx = 3523
    #10;
    addra = 32'd112768;
    dina = {96'd0, 16'd39854, 16'd56037, 16'd41223, 16'd62766, 16'd289, 16'd54779, 16'd16985, 16'd17807, 16'd4489, 16'd16990}; // indx = 3524
    #10;
    addra = 32'd112800;
    dina = {96'd0, 16'd12709, 16'd45803, 16'd21910, 16'd15804, 16'd6205, 16'd8816, 16'd63115, 16'd17398, 16'd42832, 16'd25613}; // indx = 3525
    #10;
    addra = 32'd112832;
    dina = {96'd0, 16'd54182, 16'd8468, 16'd28149, 16'd20143, 16'd479, 16'd50900, 16'd32538, 16'd49033, 16'd18464, 16'd9938}; // indx = 3526
    #10;
    addra = 32'd112864;
    dina = {96'd0, 16'd34224, 16'd19876, 16'd5226, 16'd60874, 16'd12060, 16'd25184, 16'd62727, 16'd40239, 16'd33803, 16'd42010}; // indx = 3527
    #10;
    addra = 32'd112896;
    dina = {96'd0, 16'd8532, 16'd1095, 16'd21928, 16'd58597, 16'd14596, 16'd1529, 16'd46412, 16'd19665, 16'd38717, 16'd7472}; // indx = 3528
    #10;
    addra = 32'd112928;
    dina = {96'd0, 16'd27292, 16'd643, 16'd5822, 16'd23145, 16'd36663, 16'd56808, 16'd42638, 16'd2471, 16'd7453, 16'd51741}; // indx = 3529
    #10;
    addra = 32'd112960;
    dina = {96'd0, 16'd5836, 16'd43971, 16'd63043, 16'd14686, 16'd29175, 16'd11428, 16'd49603, 16'd53019, 16'd27491, 16'd7536}; // indx = 3530
    #10;
    addra = 32'd112992;
    dina = {96'd0, 16'd44196, 16'd42775, 16'd50483, 16'd24788, 16'd49242, 16'd37294, 16'd57680, 16'd62199, 16'd60905, 16'd50757}; // indx = 3531
    #10;
    addra = 32'd113024;
    dina = {96'd0, 16'd40605, 16'd40103, 16'd53235, 16'd33272, 16'd9503, 16'd6770, 16'd369, 16'd61409, 16'd14221, 16'd49845}; // indx = 3532
    #10;
    addra = 32'd113056;
    dina = {96'd0, 16'd13816, 16'd49484, 16'd18296, 16'd101, 16'd371, 16'd4648, 16'd37328, 16'd61524, 16'd41238, 16'd20202}; // indx = 3533
    #10;
    addra = 32'd113088;
    dina = {96'd0, 16'd15219, 16'd13415, 16'd5088, 16'd20706, 16'd53023, 16'd53127, 16'd44577, 16'd28733, 16'd58688, 16'd40744}; // indx = 3534
    #10;
    addra = 32'd113120;
    dina = {96'd0, 16'd20992, 16'd31028, 16'd58567, 16'd34806, 16'd56737, 16'd51530, 16'd27299, 16'd49302, 16'd26095, 16'd28047}; // indx = 3535
    #10;
    addra = 32'd113152;
    dina = {96'd0, 16'd42195, 16'd45499, 16'd38698, 16'd12469, 16'd59502, 16'd17777, 16'd4946, 16'd56544, 16'd44412, 16'd45964}; // indx = 3536
    #10;
    addra = 32'd113184;
    dina = {96'd0, 16'd23697, 16'd36712, 16'd7250, 16'd28483, 16'd13678, 16'd10853, 16'd36118, 16'd60919, 16'd38328, 16'd26900}; // indx = 3537
    #10;
    addra = 32'd113216;
    dina = {96'd0, 16'd26327, 16'd58279, 16'd34212, 16'd48342, 16'd37737, 16'd46246, 16'd37012, 16'd33900, 16'd37186, 16'd9445}; // indx = 3538
    #10;
    addra = 32'd113248;
    dina = {96'd0, 16'd54884, 16'd19489, 16'd49698, 16'd44067, 16'd45446, 16'd9214, 16'd39585, 16'd14569, 16'd34572, 16'd20115}; // indx = 3539
    #10;
    addra = 32'd113280;
    dina = {96'd0, 16'd35570, 16'd53528, 16'd56560, 16'd30323, 16'd7441, 16'd53582, 16'd43604, 16'd23751, 16'd51695, 16'd30125}; // indx = 3540
    #10;
    addra = 32'd113312;
    dina = {96'd0, 16'd45044, 16'd51176, 16'd64201, 16'd259, 16'd41637, 16'd49744, 16'd62363, 16'd57828, 16'd24775, 16'd49248}; // indx = 3541
    #10;
    addra = 32'd113344;
    dina = {96'd0, 16'd436, 16'd32223, 16'd22066, 16'd28997, 16'd31823, 16'd20123, 16'd27665, 16'd27002, 16'd9137, 16'd19437}; // indx = 3542
    #10;
    addra = 32'd113376;
    dina = {96'd0, 16'd49671, 16'd11097, 16'd32592, 16'd31658, 16'd8812, 16'd27565, 16'd37368, 16'd37312, 16'd33430, 16'd26557}; // indx = 3543
    #10;
    addra = 32'd113408;
    dina = {96'd0, 16'd59072, 16'd46375, 16'd50554, 16'd20462, 16'd13772, 16'd57506, 16'd32493, 16'd6380, 16'd43518, 16'd7385}; // indx = 3544
    #10;
    addra = 32'd113440;
    dina = {96'd0, 16'd62417, 16'd50841, 16'd11307, 16'd60354, 16'd20361, 16'd13990, 16'd2589, 16'd18579, 16'd50939, 16'd12475}; // indx = 3545
    #10;
    addra = 32'd113472;
    dina = {96'd0, 16'd35358, 16'd45071, 16'd6098, 16'd12424, 16'd25586, 16'd43107, 16'd60661, 16'd51427, 16'd12724, 16'd52092}; // indx = 3546
    #10;
    addra = 32'd113504;
    dina = {96'd0, 16'd15029, 16'd7663, 16'd19664, 16'd46330, 16'd2364, 16'd62881, 16'd1117, 16'd48711, 16'd60146, 16'd14788}; // indx = 3547
    #10;
    addra = 32'd113536;
    dina = {96'd0, 16'd36753, 16'd39723, 16'd28939, 16'd18440, 16'd9090, 16'd25881, 16'd38451, 16'd40698, 16'd1144, 16'd23364}; // indx = 3548
    #10;
    addra = 32'd113568;
    dina = {96'd0, 16'd23910, 16'd60653, 16'd16394, 16'd42048, 16'd29072, 16'd12666, 16'd50252, 16'd36092, 16'd32795, 16'd64880}; // indx = 3549
    #10;
    addra = 32'd113600;
    dina = {96'd0, 16'd21044, 16'd53196, 16'd18933, 16'd15331, 16'd65283, 16'd57265, 16'd21012, 16'd33321, 16'd55153, 16'd53609}; // indx = 3550
    #10;
    addra = 32'd113632;
    dina = {96'd0, 16'd51430, 16'd42877, 16'd39672, 16'd8790, 16'd22099, 16'd63184, 16'd3860, 16'd27305, 16'd60868, 16'd59039}; // indx = 3551
    #10;
    addra = 32'd113664;
    dina = {96'd0, 16'd10871, 16'd27945, 16'd36986, 16'd47174, 16'd7911, 16'd16164, 16'd60979, 16'd51138, 16'd57287, 16'd27383}; // indx = 3552
    #10;
    addra = 32'd113696;
    dina = {96'd0, 16'd55272, 16'd32318, 16'd5851, 16'd61264, 16'd14007, 16'd32482, 16'd58935, 16'd21613, 16'd24255, 16'd51158}; // indx = 3553
    #10;
    addra = 32'd113728;
    dina = {96'd0, 16'd5234, 16'd20488, 16'd29144, 16'd30369, 16'd6875, 16'd32619, 16'd14346, 16'd41057, 16'd50756, 16'd938}; // indx = 3554
    #10;
    addra = 32'd113760;
    dina = {96'd0, 16'd54117, 16'd61575, 16'd47670, 16'd5876, 16'd26371, 16'd45018, 16'd22559, 16'd38662, 16'd61719, 16'd51724}; // indx = 3555
    #10;
    addra = 32'd113792;
    dina = {96'd0, 16'd30907, 16'd30698, 16'd41634, 16'd16096, 16'd54357, 16'd15688, 16'd7905, 16'd35276, 16'd16907, 16'd27432}; // indx = 3556
    #10;
    addra = 32'd113824;
    dina = {96'd0, 16'd60606, 16'd32110, 16'd58049, 16'd22633, 16'd26156, 16'd60383, 16'd34269, 16'd11030, 16'd55333, 16'd61126}; // indx = 3557
    #10;
    addra = 32'd113856;
    dina = {96'd0, 16'd12399, 16'd44931, 16'd8138, 16'd37637, 16'd57290, 16'd51806, 16'd49202, 16'd7665, 16'd33164, 16'd36730}; // indx = 3558
    #10;
    addra = 32'd113888;
    dina = {96'd0, 16'd4287, 16'd31227, 16'd40923, 16'd34560, 16'd44896, 16'd21984, 16'd34907, 16'd14139, 16'd174, 16'd21461}; // indx = 3559
    #10;
    addra = 32'd113920;
    dina = {96'd0, 16'd52183, 16'd59484, 16'd17198, 16'd42923, 16'd55021, 16'd4130, 16'd25617, 16'd45236, 16'd41176, 16'd62617}; // indx = 3560
    #10;
    addra = 32'd113952;
    dina = {96'd0, 16'd5922, 16'd62454, 16'd1120, 16'd20656, 16'd60889, 16'd56297, 16'd42881, 16'd58704, 16'd31839, 16'd25822}; // indx = 3561
    #10;
    addra = 32'd113984;
    dina = {96'd0, 16'd60695, 16'd44111, 16'd21530, 16'd49117, 16'd50991, 16'd31319, 16'd10275, 16'd37417, 16'd56294, 16'd13694}; // indx = 3562
    #10;
    addra = 32'd114016;
    dina = {96'd0, 16'd28954, 16'd22267, 16'd24574, 16'd62517, 16'd33011, 16'd39846, 16'd16636, 16'd40374, 16'd39939, 16'd9724}; // indx = 3563
    #10;
    addra = 32'd114048;
    dina = {96'd0, 16'd5637, 16'd19359, 16'd14932, 16'd10827, 16'd41812, 16'd62407, 16'd35920, 16'd8507, 16'd6664, 16'd64267}; // indx = 3564
    #10;
    addra = 32'd114080;
    dina = {96'd0, 16'd41035, 16'd1166, 16'd48651, 16'd25022, 16'd63602, 16'd26757, 16'd44817, 16'd39414, 16'd46430, 16'd1866}; // indx = 3565
    #10;
    addra = 32'd114112;
    dina = {96'd0, 16'd3624, 16'd34142, 16'd37940, 16'd49766, 16'd37836, 16'd31989, 16'd42978, 16'd8748, 16'd46241, 16'd42374}; // indx = 3566
    #10;
    addra = 32'd114144;
    dina = {96'd0, 16'd15488, 16'd21923, 16'd41541, 16'd22056, 16'd55386, 16'd23086, 16'd28194, 16'd6311, 16'd46560, 16'd48633}; // indx = 3567
    #10;
    addra = 32'd114176;
    dina = {96'd0, 16'd23102, 16'd20888, 16'd26940, 16'd10857, 16'd52033, 16'd731, 16'd34701, 16'd25855, 16'd55457, 16'd12516}; // indx = 3568
    #10;
    addra = 32'd114208;
    dina = {96'd0, 16'd55641, 16'd33998, 16'd11535, 16'd34526, 16'd43961, 16'd1991, 16'd39590, 16'd53837, 16'd59051, 16'd22360}; // indx = 3569
    #10;
    addra = 32'd114240;
    dina = {96'd0, 16'd2373, 16'd64193, 16'd54952, 16'd10211, 16'd30529, 16'd22205, 16'd62236, 16'd49479, 16'd10350, 16'd27766}; // indx = 3570
    #10;
    addra = 32'd114272;
    dina = {96'd0, 16'd35632, 16'd33979, 16'd27753, 16'd40646, 16'd40666, 16'd21981, 16'd32440, 16'd54190, 16'd46577, 16'd47729}; // indx = 3571
    #10;
    addra = 32'd114304;
    dina = {96'd0, 16'd36205, 16'd14594, 16'd15063, 16'd39290, 16'd63693, 16'd59091, 16'd59335, 16'd14659, 16'd13856, 16'd3620}; // indx = 3572
    #10;
    addra = 32'd114336;
    dina = {96'd0, 16'd47622, 16'd10963, 16'd15275, 16'd18430, 16'd23489, 16'd13339, 16'd28940, 16'd27396, 16'd27007, 16'd46903}; // indx = 3573
    #10;
    addra = 32'd114368;
    dina = {96'd0, 16'd12395, 16'd60837, 16'd26450, 16'd32121, 16'd61370, 16'd31265, 16'd52980, 16'd54939, 16'd34540, 16'd29116}; // indx = 3574
    #10;
    addra = 32'd114400;
    dina = {96'd0, 16'd20882, 16'd16824, 16'd47078, 16'd3320, 16'd12515, 16'd698, 16'd25534, 16'd31431, 16'd46510, 16'd11870}; // indx = 3575
    #10;
    addra = 32'd114432;
    dina = {96'd0, 16'd49963, 16'd62016, 16'd44021, 16'd22491, 16'd56117, 16'd15491, 16'd28477, 16'd47478, 16'd3197, 16'd60813}; // indx = 3576
    #10;
    addra = 32'd114464;
    dina = {96'd0, 16'd38411, 16'd33345, 16'd62428, 16'd9147, 16'd32337, 16'd49668, 16'd40724, 16'd37176, 16'd63652, 16'd64750}; // indx = 3577
    #10;
    addra = 32'd114496;
    dina = {96'd0, 16'd51591, 16'd16128, 16'd4808, 16'd48044, 16'd35058, 16'd60946, 16'd64819, 16'd42261, 16'd29844, 16'd51513}; // indx = 3578
    #10;
    addra = 32'd114528;
    dina = {96'd0, 16'd61247, 16'd63207, 16'd1158, 16'd38416, 16'd47506, 16'd4586, 16'd39970, 16'd14833, 16'd4136, 16'd35332}; // indx = 3579
    #10;
    addra = 32'd114560;
    dina = {96'd0, 16'd36130, 16'd49549, 16'd18661, 16'd18634, 16'd4432, 16'd6435, 16'd8996, 16'd22952, 16'd23755, 16'd62380}; // indx = 3580
    #10;
    addra = 32'd114592;
    dina = {96'd0, 16'd21566, 16'd63757, 16'd10692, 16'd27380, 16'd25291, 16'd47580, 16'd63564, 16'd25199, 16'd64507, 16'd39404}; // indx = 3581
    #10;
    addra = 32'd114624;
    dina = {96'd0, 16'd42361, 16'd41726, 16'd64096, 16'd63913, 16'd59040, 16'd43823, 16'd20508, 16'd10800, 16'd32993, 16'd9960}; // indx = 3582
    #10;
    addra = 32'd114656;
    dina = {96'd0, 16'd61837, 16'd31441, 16'd53244, 16'd24920, 16'd20575, 16'd46930, 16'd10722, 16'd28870, 16'd43249, 16'd52718}; // indx = 3583
    #10;
    addra = 32'd114688;
    dina = {96'd0, 16'd14652, 16'd15155, 16'd53614, 16'd49242, 16'd20415, 16'd3866, 16'd31980, 16'd17147, 16'd27450, 16'd51575}; // indx = 3584
    #10;
    addra = 32'd114720;
    dina = {96'd0, 16'd20357, 16'd56711, 16'd54836, 16'd17052, 16'd54415, 16'd63352, 16'd58285, 16'd20349, 16'd28702, 16'd34976}; // indx = 3585
    #10;
    addra = 32'd114752;
    dina = {96'd0, 16'd20789, 16'd47500, 16'd64410, 16'd40797, 16'd17529, 16'd44691, 16'd7357, 16'd62797, 16'd7666, 16'd3265}; // indx = 3586
    #10;
    addra = 32'd114784;
    dina = {96'd0, 16'd35631, 16'd44790, 16'd30298, 16'd45473, 16'd14100, 16'd124, 16'd42222, 16'd7593, 16'd44201, 16'd54090}; // indx = 3587
    #10;
    addra = 32'd114816;
    dina = {96'd0, 16'd37063, 16'd31935, 16'd50655, 16'd21769, 16'd36642, 16'd21351, 16'd42813, 16'd10836, 16'd38824, 16'd27891}; // indx = 3588
    #10;
    addra = 32'd114848;
    dina = {96'd0, 16'd43084, 16'd45915, 16'd51828, 16'd34493, 16'd42328, 16'd15774, 16'd4270, 16'd38390, 16'd37379, 16'd2214}; // indx = 3589
    #10;
    addra = 32'd114880;
    dina = {96'd0, 16'd27066, 16'd16352, 16'd469, 16'd23683, 16'd40391, 16'd51740, 16'd41229, 16'd29126, 16'd9906, 16'd5243}; // indx = 3590
    #10;
    addra = 32'd114912;
    dina = {96'd0, 16'd63203, 16'd49234, 16'd12409, 16'd24517, 16'd65433, 16'd1209, 16'd7966, 16'd30603, 16'd5428, 16'd27516}; // indx = 3591
    #10;
    addra = 32'd114944;
    dina = {96'd0, 16'd59103, 16'd64364, 16'd5670, 16'd39437, 16'd37658, 16'd57113, 16'd35879, 16'd1108, 16'd23573, 16'd62478}; // indx = 3592
    #10;
    addra = 32'd114976;
    dina = {96'd0, 16'd12178, 16'd28076, 16'd9999, 16'd27723, 16'd23333, 16'd18295, 16'd10988, 16'd15376, 16'd2808, 16'd10969}; // indx = 3593
    #10;
    addra = 32'd115008;
    dina = {96'd0, 16'd8951, 16'd34050, 16'd15809, 16'd9439, 16'd50415, 16'd17299, 16'd40420, 16'd43888, 16'd59408, 16'd40097}; // indx = 3594
    #10;
    addra = 32'd115040;
    dina = {96'd0, 16'd12330, 16'd15629, 16'd27655, 16'd39592, 16'd36274, 16'd37962, 16'd9728, 16'd34256, 16'd4716, 16'd57370}; // indx = 3595
    #10;
    addra = 32'd115072;
    dina = {96'd0, 16'd65454, 16'd16830, 16'd61341, 16'd308, 16'd62068, 16'd30848, 16'd59677, 16'd48299, 16'd56223, 16'd53641}; // indx = 3596
    #10;
    addra = 32'd115104;
    dina = {96'd0, 16'd26396, 16'd3871, 16'd18250, 16'd8354, 16'd34989, 16'd28004, 16'd3533, 16'd9241, 16'd63519, 16'd20050}; // indx = 3597
    #10;
    addra = 32'd115136;
    dina = {96'd0, 16'd3494, 16'd20364, 16'd11599, 16'd58340, 16'd53616, 16'd27493, 16'd32636, 16'd16792, 16'd9594, 16'd3063}; // indx = 3598
    #10;
    addra = 32'd115168;
    dina = {96'd0, 16'd13398, 16'd7718, 16'd35069, 16'd44659, 16'd20931, 16'd62579, 16'd38063, 16'd57838, 16'd42962, 16'd22102}; // indx = 3599
    #10;
    addra = 32'd115200;
    dina = {96'd0, 16'd64763, 16'd3993, 16'd32058, 16'd20722, 16'd65013, 16'd53257, 16'd28825, 16'd23914, 16'd42147, 16'd43549}; // indx = 3600
    #10;
    addra = 32'd115232;
    dina = {96'd0, 16'd34131, 16'd13578, 16'd60040, 16'd56232, 16'd48675, 16'd63745, 16'd49290, 16'd17832, 16'd6881, 16'd29252}; // indx = 3601
    #10;
    addra = 32'd115264;
    dina = {96'd0, 16'd20100, 16'd64098, 16'd30072, 16'd86, 16'd30118, 16'd38615, 16'd11391, 16'd37818, 16'd63613, 16'd51742}; // indx = 3602
    #10;
    addra = 32'd115296;
    dina = {96'd0, 16'd10738, 16'd15604, 16'd17977, 16'd22290, 16'd56025, 16'd34540, 16'd26528, 16'd42341, 16'd62052, 16'd33051}; // indx = 3603
    #10;
    addra = 32'd115328;
    dina = {96'd0, 16'd50855, 16'd53366, 16'd33297, 16'd2689, 16'd19265, 16'd22601, 16'd38113, 16'd8151, 16'd37534, 16'd38525}; // indx = 3604
    #10;
    addra = 32'd115360;
    dina = {96'd0, 16'd57108, 16'd56719, 16'd40467, 16'd5479, 16'd24552, 16'd30899, 16'd61563, 16'd44321, 16'd52375, 16'd33031}; // indx = 3605
    #10;
    addra = 32'd115392;
    dina = {96'd0, 16'd25668, 16'd17430, 16'd8604, 16'd17916, 16'd42235, 16'd8734, 16'd13, 16'd2229, 16'd10600, 16'd50283}; // indx = 3606
    #10;
    addra = 32'd115424;
    dina = {96'd0, 16'd26033, 16'd17934, 16'd51223, 16'd15092, 16'd48812, 16'd48160, 16'd4323, 16'd10629, 16'd38301, 16'd61558}; // indx = 3607
    #10;
    addra = 32'd115456;
    dina = {96'd0, 16'd22864, 16'd53497, 16'd36229, 16'd40051, 16'd52160, 16'd45617, 16'd59380, 16'd50532, 16'd6196, 16'd18531}; // indx = 3608
    #10;
    addra = 32'd115488;
    dina = {96'd0, 16'd4786, 16'd27021, 16'd5722, 16'd16023, 16'd43944, 16'd40951, 16'd43416, 16'd13712, 16'd35141, 16'd55772}; // indx = 3609
    #10;
    addra = 32'd115520;
    dina = {96'd0, 16'd19699, 16'd60824, 16'd23596, 16'd43985, 16'd44663, 16'd29137, 16'd50649, 16'd44607, 16'd36661, 16'd26412}; // indx = 3610
    #10;
    addra = 32'd115552;
    dina = {96'd0, 16'd33464, 16'd15437, 16'd54940, 16'd7531, 16'd12160, 16'd43019, 16'd25774, 16'd6450, 16'd64497, 16'd56456}; // indx = 3611
    #10;
    addra = 32'd115584;
    dina = {96'd0, 16'd30969, 16'd42058, 16'd54945, 16'd54762, 16'd26336, 16'd10918, 16'd40675, 16'd59004, 16'd40301, 16'd53525}; // indx = 3612
    #10;
    addra = 32'd115616;
    dina = {96'd0, 16'd5568, 16'd61163, 16'd42717, 16'd21636, 16'd6088, 16'd2893, 16'd41201, 16'd65002, 16'd26001, 16'd4450}; // indx = 3613
    #10;
    addra = 32'd115648;
    dina = {96'd0, 16'd14733, 16'd9237, 16'd13566, 16'd43787, 16'd17144, 16'd13561, 16'd17747, 16'd15538, 16'd25718, 16'd37629}; // indx = 3614
    #10;
    addra = 32'd115680;
    dina = {96'd0, 16'd48737, 16'd26440, 16'd50000, 16'd50808, 16'd62388, 16'd49210, 16'd5117, 16'd30061, 16'd65425, 16'd33137}; // indx = 3615
    #10;
    addra = 32'd115712;
    dina = {96'd0, 16'd62956, 16'd60199, 16'd2097, 16'd28370, 16'd47886, 16'd6599, 16'd53956, 16'd9770, 16'd4479, 16'd62713}; // indx = 3616
    #10;
    addra = 32'd115744;
    dina = {96'd0, 16'd29367, 16'd57601, 16'd30825, 16'd27511, 16'd52375, 16'd18597, 16'd45118, 16'd36056, 16'd18247, 16'd37962}; // indx = 3617
    #10;
    addra = 32'd115776;
    dina = {96'd0, 16'd8605, 16'd5388, 16'd61700, 16'd32130, 16'd16130, 16'd17755, 16'd56758, 16'd46798, 16'd39175, 16'd7894}; // indx = 3618
    #10;
    addra = 32'd115808;
    dina = {96'd0, 16'd54694, 16'd12197, 16'd54058, 16'd52487, 16'd3190, 16'd11359, 16'd56496, 16'd63540, 16'd63713, 16'd15597}; // indx = 3619
    #10;
    addra = 32'd115840;
    dina = {96'd0, 16'd35590, 16'd657, 16'd39456, 16'd51047, 16'd31223, 16'd45350, 16'd6124, 16'd24750, 16'd9415, 16'd46100}; // indx = 3620
    #10;
    addra = 32'd115872;
    dina = {96'd0, 16'd32417, 16'd43936, 16'd23994, 16'd41993, 16'd48398, 16'd51249, 16'd49578, 16'd5850, 16'd49913, 16'd47742}; // indx = 3621
    #10;
    addra = 32'd115904;
    dina = {96'd0, 16'd30066, 16'd52654, 16'd35900, 16'd19664, 16'd62629, 16'd22144, 16'd33833, 16'd27239, 16'd23190, 16'd63855}; // indx = 3622
    #10;
    addra = 32'd115936;
    dina = {96'd0, 16'd36468, 16'd19314, 16'd20710, 16'd23518, 16'd13830, 16'd5596, 16'd35424, 16'd33023, 16'd21697, 16'd54729}; // indx = 3623
    #10;
    addra = 32'd115968;
    dina = {96'd0, 16'd3798, 16'd18241, 16'd13306, 16'd39180, 16'd38507, 16'd18547, 16'd39118, 16'd33693, 16'd34300, 16'd49668}; // indx = 3624
    #10;
    addra = 32'd116000;
    dina = {96'd0, 16'd61338, 16'd39173, 16'd27696, 16'd1732, 16'd64513, 16'd13425, 16'd39208, 16'd29099, 16'd60369, 16'd22166}; // indx = 3625
    #10;
    addra = 32'd116032;
    dina = {96'd0, 16'd65441, 16'd48864, 16'd27249, 16'd31876, 16'd63093, 16'd8096, 16'd18153, 16'd2641, 16'd15561, 16'd5977}; // indx = 3626
    #10;
    addra = 32'd116064;
    dina = {96'd0, 16'd50698, 16'd30732, 16'd13540, 16'd12854, 16'd38265, 16'd3293, 16'd20260, 16'd6416, 16'd27502, 16'd28322}; // indx = 3627
    #10;
    addra = 32'd116096;
    dina = {96'd0, 16'd20449, 16'd528, 16'd45385, 16'd56689, 16'd10677, 16'd48698, 16'd16367, 16'd29381, 16'd21728, 16'd35997}; // indx = 3628
    #10;
    addra = 32'd116128;
    dina = {96'd0, 16'd35899, 16'd15205, 16'd13915, 16'd10342, 16'd12849, 16'd4587, 16'd21020, 16'd33375, 16'd27396, 16'd53043}; // indx = 3629
    #10;
    addra = 32'd116160;
    dina = {96'd0, 16'd23726, 16'd23436, 16'd64283, 16'd28837, 16'd31505, 16'd15005, 16'd28720, 16'd60189, 16'd3222, 16'd1592}; // indx = 3630
    #10;
    addra = 32'd116192;
    dina = {96'd0, 16'd22194, 16'd49129, 16'd34752, 16'd7543, 16'd4791, 16'd42884, 16'd17002, 16'd30765, 16'd18899, 16'd60010}; // indx = 3631
    #10;
    addra = 32'd116224;
    dina = {96'd0, 16'd35296, 16'd18021, 16'd54372, 16'd32652, 16'd17764, 16'd23176, 16'd50500, 16'd40475, 16'd10572, 16'd2827}; // indx = 3632
    #10;
    addra = 32'd116256;
    dina = {96'd0, 16'd13265, 16'd38500, 16'd39790, 16'd50272, 16'd4062, 16'd21421, 16'd28944, 16'd35850, 16'd3078, 16'd11023}; // indx = 3633
    #10;
    addra = 32'd116288;
    dina = {96'd0, 16'd63403, 16'd48042, 16'd50479, 16'd39303, 16'd47150, 16'd35659, 16'd16265, 16'd59177, 16'd54718, 16'd39590}; // indx = 3634
    #10;
    addra = 32'd116320;
    dina = {96'd0, 16'd7435, 16'd42196, 16'd50533, 16'd62637, 16'd63318, 16'd7386, 16'd32747, 16'd46815, 16'd41731, 16'd49692}; // indx = 3635
    #10;
    addra = 32'd116352;
    dina = {96'd0, 16'd59797, 16'd3328, 16'd64233, 16'd33641, 16'd50414, 16'd32768, 16'd52122, 16'd5595, 16'd54716, 16'd48441}; // indx = 3636
    #10;
    addra = 32'd116384;
    dina = {96'd0, 16'd38018, 16'd666, 16'd31750, 16'd39126, 16'd60835, 16'd45147, 16'd57428, 16'd37945, 16'd9665, 16'd16292}; // indx = 3637
    #10;
    addra = 32'd116416;
    dina = {96'd0, 16'd50676, 16'd15686, 16'd19329, 16'd14839, 16'd53775, 16'd54665, 16'd60238, 16'd36126, 16'd27873, 16'd62204}; // indx = 3638
    #10;
    addra = 32'd116448;
    dina = {96'd0, 16'd20798, 16'd18640, 16'd10911, 16'd19536, 16'd25303, 16'd34454, 16'd16053, 16'd53784, 16'd48514, 16'd8791}; // indx = 3639
    #10;
    addra = 32'd116480;
    dina = {96'd0, 16'd45358, 16'd22623, 16'd37211, 16'd55003, 16'd61384, 16'd16725, 16'd26812, 16'd46940, 16'd31841, 16'd53372}; // indx = 3640
    #10;
    addra = 32'd116512;
    dina = {96'd0, 16'd42927, 16'd31084, 16'd36938, 16'd45629, 16'd13357, 16'd46353, 16'd1246, 16'd51655, 16'd37734, 16'd52885}; // indx = 3641
    #10;
    addra = 32'd116544;
    dina = {96'd0, 16'd48211, 16'd43643, 16'd5671, 16'd14229, 16'd36735, 16'd36500, 16'd50798, 16'd24191, 16'd27064, 16'd56800}; // indx = 3642
    #10;
    addra = 32'd116576;
    dina = {96'd0, 16'd59657, 16'd64552, 16'd24837, 16'd45419, 16'd31191, 16'd36474, 16'd48777, 16'd12771, 16'd39354, 16'd34257}; // indx = 3643
    #10;
    addra = 32'd116608;
    dina = {96'd0, 16'd51164, 16'd63892, 16'd25719, 16'd39791, 16'd48210, 16'd4675, 16'd31989, 16'd59757, 16'd38595, 16'd24426}; // indx = 3644
    #10;
    addra = 32'd116640;
    dina = {96'd0, 16'd24105, 16'd26697, 16'd26782, 16'd63625, 16'd53197, 16'd50566, 16'd2958, 16'd54207, 16'd40822, 16'd32390}; // indx = 3645
    #10;
    addra = 32'd116672;
    dina = {96'd0, 16'd25829, 16'd57449, 16'd14261, 16'd62084, 16'd23649, 16'd34642, 16'd42677, 16'd17520, 16'd59542, 16'd28590}; // indx = 3646
    #10;
    addra = 32'd116704;
    dina = {96'd0, 16'd41804, 16'd38284, 16'd5189, 16'd48179, 16'd19694, 16'd45112, 16'd33146, 16'd34215, 16'd36552, 16'd57839}; // indx = 3647
    #10;
    addra = 32'd116736;
    dina = {96'd0, 16'd29263, 16'd56705, 16'd25731, 16'd5089, 16'd22878, 16'd63677, 16'd30583, 16'd57457, 16'd30796, 16'd43049}; // indx = 3648
    #10;
    addra = 32'd116768;
    dina = {96'd0, 16'd58869, 16'd2000, 16'd16602, 16'd34201, 16'd46482, 16'd14322, 16'd56559, 16'd60532, 16'd2455, 16'd34980}; // indx = 3649
    #10;
    addra = 32'd116800;
    dina = {96'd0, 16'd50590, 16'd30503, 16'd3072, 16'd43614, 16'd22333, 16'd56823, 16'd11637, 16'd57533, 16'd39099, 16'd28464}; // indx = 3650
    #10;
    addra = 32'd116832;
    dina = {96'd0, 16'd25469, 16'd37693, 16'd34825, 16'd38860, 16'd41411, 16'd11226, 16'd56178, 16'd30024, 16'd10634, 16'd49175}; // indx = 3651
    #10;
    addra = 32'd116864;
    dina = {96'd0, 16'd17229, 16'd53186, 16'd45536, 16'd40293, 16'd42556, 16'd24494, 16'd17227, 16'd42312, 16'd51649, 16'd13998}; // indx = 3652
    #10;
    addra = 32'd116896;
    dina = {96'd0, 16'd61257, 16'd5295, 16'd26426, 16'd42467, 16'd8926, 16'd2571, 16'd37929, 16'd11253, 16'd867, 16'd52110}; // indx = 3653
    #10;
    addra = 32'd116928;
    dina = {96'd0, 16'd58669, 16'd61213, 16'd16051, 16'd86, 16'd36130, 16'd47620, 16'd43318, 16'd12444, 16'd39252, 16'd43101}; // indx = 3654
    #10;
    addra = 32'd116960;
    dina = {96'd0, 16'd58268, 16'd4656, 16'd26601, 16'd36710, 16'd62024, 16'd37919, 16'd44539, 16'd19986, 16'd23180, 16'd62889}; // indx = 3655
    #10;
    addra = 32'd116992;
    dina = {96'd0, 16'd33880, 16'd45555, 16'd23929, 16'd20455, 16'd44392, 16'd18984, 16'd9653, 16'd57995, 16'd58875, 16'd49820}; // indx = 3656
    #10;
    addra = 32'd117024;
    dina = {96'd0, 16'd52356, 16'd20895, 16'd12518, 16'd30158, 16'd31761, 16'd38936, 16'd46231, 16'd13337, 16'd60121, 16'd12643}; // indx = 3657
    #10;
    addra = 32'd117056;
    dina = {96'd0, 16'd26655, 16'd59545, 16'd22839, 16'd22766, 16'd52281, 16'd46224, 16'd39189, 16'd3848, 16'd19676, 16'd26575}; // indx = 3658
    #10;
    addra = 32'd117088;
    dina = {96'd0, 16'd27161, 16'd21542, 16'd56727, 16'd52272, 16'd48255, 16'd11031, 16'd43698, 16'd63135, 16'd54759, 16'd10918}; // indx = 3659
    #10;
    addra = 32'd117120;
    dina = {96'd0, 16'd57375, 16'd6675, 16'd15424, 16'd27149, 16'd32828, 16'd58673, 16'd5454, 16'd51042, 16'd45821, 16'd36709}; // indx = 3660
    #10;
    addra = 32'd117152;
    dina = {96'd0, 16'd50811, 16'd5607, 16'd59051, 16'd59636, 16'd59475, 16'd50030, 16'd50222, 16'd24635, 16'd28490, 16'd49102}; // indx = 3661
    #10;
    addra = 32'd117184;
    dina = {96'd0, 16'd10610, 16'd9101, 16'd32479, 16'd4220, 16'd8352, 16'd34321, 16'd64904, 16'd52910, 16'd57527, 16'd26341}; // indx = 3662
    #10;
    addra = 32'd117216;
    dina = {96'd0, 16'd44882, 16'd64546, 16'd8200, 16'd44623, 16'd38070, 16'd8723, 16'd4453, 16'd65210, 16'd40682, 16'd32844}; // indx = 3663
    #10;
    addra = 32'd117248;
    dina = {96'd0, 16'd26902, 16'd43171, 16'd16365, 16'd37419, 16'd65226, 16'd3003, 16'd51200, 16'd2842, 16'd55401, 16'd32321}; // indx = 3664
    #10;
    addra = 32'd117280;
    dina = {96'd0, 16'd46430, 16'd49653, 16'd23433, 16'd50007, 16'd25694, 16'd8067, 16'd21787, 16'd38566, 16'd5280, 16'd27108}; // indx = 3665
    #10;
    addra = 32'd117312;
    dina = {96'd0, 16'd44573, 16'd59186, 16'd53827, 16'd64767, 16'd18243, 16'd6984, 16'd50989, 16'd9348, 16'd21844, 16'd22851}; // indx = 3666
    #10;
    addra = 32'd117344;
    dina = {96'd0, 16'd55807, 16'd50218, 16'd23673, 16'd30608, 16'd56166, 16'd6498, 16'd45245, 16'd30983, 16'd2631, 16'd42355}; // indx = 3667
    #10;
    addra = 32'd117376;
    dina = {96'd0, 16'd20109, 16'd37148, 16'd8539, 16'd8333, 16'd8039, 16'd37459, 16'd43108, 16'd36091, 16'd13483, 16'd49377}; // indx = 3668
    #10;
    addra = 32'd117408;
    dina = {96'd0, 16'd55201, 16'd60937, 16'd32204, 16'd9221, 16'd39118, 16'd53747, 16'd11509, 16'd26618, 16'd57263, 16'd54824}; // indx = 3669
    #10;
    addra = 32'd117440;
    dina = {96'd0, 16'd22047, 16'd60531, 16'd65533, 16'd47509, 16'd18550, 16'd65288, 16'd40348, 16'd11570, 16'd17358, 16'd44384}; // indx = 3670
    #10;
    addra = 32'd117472;
    dina = {96'd0, 16'd61222, 16'd13606, 16'd64342, 16'd7207, 16'd55907, 16'd16616, 16'd15745, 16'd9515, 16'd12129, 16'd53794}; // indx = 3671
    #10;
    addra = 32'd117504;
    dina = {96'd0, 16'd56277, 16'd60878, 16'd12069, 16'd52158, 16'd4329, 16'd44773, 16'd14061, 16'd5705, 16'd62504, 16'd21012}; // indx = 3672
    #10;
    addra = 32'd117536;
    dina = {96'd0, 16'd41363, 16'd47814, 16'd28311, 16'd20675, 16'd25916, 16'd41410, 16'd50008, 16'd50246, 16'd49115, 16'd21774}; // indx = 3673
    #10;
    addra = 32'd117568;
    dina = {96'd0, 16'd24415, 16'd52887, 16'd12377, 16'd48162, 16'd24175, 16'd11818, 16'd28687, 16'd23117, 16'd4514, 16'd3526}; // indx = 3674
    #10;
    addra = 32'd117600;
    dina = {96'd0, 16'd62216, 16'd45271, 16'd13552, 16'd26555, 16'd57873, 16'd61480, 16'd1613, 16'd13812, 16'd30653, 16'd39596}; // indx = 3675
    #10;
    addra = 32'd117632;
    dina = {96'd0, 16'd15448, 16'd43200, 16'd65149, 16'd41487, 16'd24471, 16'd25387, 16'd49520, 16'd30580, 16'd6267, 16'd2032}; // indx = 3676
    #10;
    addra = 32'd117664;
    dina = {96'd0, 16'd51387, 16'd58892, 16'd36449, 16'd17693, 16'd52992, 16'd6104, 16'd62935, 16'd50944, 16'd24965, 16'd9781}; // indx = 3677
    #10;
    addra = 32'd117696;
    dina = {96'd0, 16'd64328, 16'd22420, 16'd13274, 16'd15372, 16'd1773, 16'd41732, 16'd5289, 16'd24842, 16'd48218, 16'd61648}; // indx = 3678
    #10;
    addra = 32'd117728;
    dina = {96'd0, 16'd59235, 16'd33279, 16'd49965, 16'd26051, 16'd6525, 16'd38480, 16'd25249, 16'd15001, 16'd57472, 16'd19066}; // indx = 3679
    #10;
    addra = 32'd117760;
    dina = {96'd0, 16'd39729, 16'd29311, 16'd29731, 16'd54761, 16'd161, 16'd21681, 16'd9673, 16'd38934, 16'd5609, 16'd39262}; // indx = 3680
    #10;
    addra = 32'd117792;
    dina = {96'd0, 16'd33997, 16'd11096, 16'd50782, 16'd27483, 16'd60437, 16'd45150, 16'd5169, 16'd62356, 16'd65400, 16'd31212}; // indx = 3681
    #10;
    addra = 32'd117824;
    dina = {96'd0, 16'd7429, 16'd10058, 16'd59868, 16'd55098, 16'd28997, 16'd51190, 16'd47808, 16'd61832, 16'd53792, 16'd58054}; // indx = 3682
    #10;
    addra = 32'd117856;
    dina = {96'd0, 16'd30302, 16'd19993, 16'd17728, 16'd54406, 16'd12663, 16'd63142, 16'd25482, 16'd22213, 16'd57686, 16'd25744}; // indx = 3683
    #10;
    addra = 32'd117888;
    dina = {96'd0, 16'd5979, 16'd35188, 16'd14717, 16'd10887, 16'd50089, 16'd24140, 16'd41303, 16'd12194, 16'd11, 16'd21563}; // indx = 3684
    #10;
    addra = 32'd117920;
    dina = {96'd0, 16'd7283, 16'd64829, 16'd32122, 16'd44830, 16'd3688, 16'd41348, 16'd22816, 16'd56939, 16'd2043, 16'd5574}; // indx = 3685
    #10;
    addra = 32'd117952;
    dina = {96'd0, 16'd20755, 16'd19700, 16'd48385, 16'd29845, 16'd47197, 16'd65131, 16'd48454, 16'd16016, 16'd20974, 16'd43324}; // indx = 3686
    #10;
    addra = 32'd117984;
    dina = {96'd0, 16'd61487, 16'd3499, 16'd21402, 16'd24365, 16'd15048, 16'd109, 16'd25024, 16'd59707, 16'd25870, 16'd19720}; // indx = 3687
    #10;
    addra = 32'd118016;
    dina = {96'd0, 16'd18459, 16'd2610, 16'd47093, 16'd10524, 16'd38100, 16'd23770, 16'd9381, 16'd33632, 16'd25626, 16'd35976}; // indx = 3688
    #10;
    addra = 32'd118048;
    dina = {96'd0, 16'd56789, 16'd61706, 16'd9883, 16'd22030, 16'd8107, 16'd63070, 16'd16831, 16'd37621, 16'd61790, 16'd49439}; // indx = 3689
    #10;
    addra = 32'd118080;
    dina = {96'd0, 16'd30556, 16'd48337, 16'd23165, 16'd41959, 16'd37763, 16'd28712, 16'd9370, 16'd46304, 16'd1096, 16'd63710}; // indx = 3690
    #10;
    addra = 32'd118112;
    dina = {96'd0, 16'd27920, 16'd54875, 16'd4838, 16'd19889, 16'd54921, 16'd40870, 16'd26668, 16'd30152, 16'd35750, 16'd39278}; // indx = 3691
    #10;
    addra = 32'd118144;
    dina = {96'd0, 16'd28331, 16'd17469, 16'd26810, 16'd21693, 16'd63547, 16'd40598, 16'd22650, 16'd4669, 16'd16891, 16'd20845}; // indx = 3692
    #10;
    addra = 32'd118176;
    dina = {96'd0, 16'd61001, 16'd33552, 16'd54582, 16'd23757, 16'd44736, 16'd22302, 16'd6550, 16'd60944, 16'd50885, 16'd183}; // indx = 3693
    #10;
    addra = 32'd118208;
    dina = {96'd0, 16'd1365, 16'd56626, 16'd49330, 16'd836, 16'd47880, 16'd7486, 16'd21161, 16'd7188, 16'd6251, 16'd37981}; // indx = 3694
    #10;
    addra = 32'd118240;
    dina = {96'd0, 16'd46183, 16'd49922, 16'd19385, 16'd58002, 16'd54060, 16'd12364, 16'd32871, 16'd12215, 16'd19677, 16'd39823}; // indx = 3695
    #10;
    addra = 32'd118272;
    dina = {96'd0, 16'd39663, 16'd45269, 16'd49145, 16'd26900, 16'd17616, 16'd33143, 16'd15476, 16'd29997, 16'd27218, 16'd59585}; // indx = 3696
    #10;
    addra = 32'd118304;
    dina = {96'd0, 16'd57925, 16'd64012, 16'd55142, 16'd14972, 16'd13895, 16'd26215, 16'd38261, 16'd50578, 16'd62710, 16'd29262}; // indx = 3697
    #10;
    addra = 32'd118336;
    dina = {96'd0, 16'd1185, 16'd4457, 16'd47179, 16'd9811, 16'd11116, 16'd6816, 16'd28015, 16'd61425, 16'd653, 16'd18140}; // indx = 3698
    #10;
    addra = 32'd118368;
    dina = {96'd0, 16'd21344, 16'd45985, 16'd13108, 16'd6839, 16'd12662, 16'd52537, 16'd57374, 16'd55621, 16'd41433, 16'd5825}; // indx = 3699
    #10;
    addra = 32'd118400;
    dina = {96'd0, 16'd18130, 16'd10477, 16'd16716, 16'd10220, 16'd61381, 16'd59294, 16'd58414, 16'd1481, 16'd16770, 16'd59583}; // indx = 3700
    #10;
    addra = 32'd118432;
    dina = {96'd0, 16'd44222, 16'd44520, 16'd19542, 16'd33594, 16'd49510, 16'd22440, 16'd32414, 16'd24511, 16'd22760, 16'd3698}; // indx = 3701
    #10;
    addra = 32'd118464;
    dina = {96'd0, 16'd43379, 16'd40037, 16'd2172, 16'd58592, 16'd47352, 16'd53214, 16'd59246, 16'd62014, 16'd55877, 16'd25061}; // indx = 3702
    #10;
    addra = 32'd118496;
    dina = {96'd0, 16'd31564, 16'd15930, 16'd60165, 16'd62342, 16'd63274, 16'd37569, 16'd36889, 16'd16557, 16'd42765, 16'd58651}; // indx = 3703
    #10;
    addra = 32'd118528;
    dina = {96'd0, 16'd56844, 16'd39873, 16'd55730, 16'd33831, 16'd42188, 16'd30810, 16'd19356, 16'd8195, 16'd13770, 16'd42858}; // indx = 3704
    #10;
    addra = 32'd118560;
    dina = {96'd0, 16'd41094, 16'd1994, 16'd65106, 16'd51335, 16'd49, 16'd41849, 16'd5054, 16'd39882, 16'd28493, 16'd64056}; // indx = 3705
    #10;
    addra = 32'd118592;
    dina = {96'd0, 16'd53979, 16'd19713, 16'd35416, 16'd16334, 16'd4647, 16'd23827, 16'd65250, 16'd54284, 16'd6191, 16'd28456}; // indx = 3706
    #10;
    addra = 32'd118624;
    dina = {96'd0, 16'd553, 16'd52168, 16'd61871, 16'd10572, 16'd17342, 16'd41249, 16'd16973, 16'd14818, 16'd38834, 16'd12858}; // indx = 3707
    #10;
    addra = 32'd118656;
    dina = {96'd0, 16'd56416, 16'd2337, 16'd35502, 16'd44564, 16'd34397, 16'd53201, 16'd19903, 16'd4825, 16'd5166, 16'd39801}; // indx = 3708
    #10;
    addra = 32'd118688;
    dina = {96'd0, 16'd24984, 16'd15292, 16'd47217, 16'd46237, 16'd13315, 16'd53091, 16'd18281, 16'd36922, 16'd35354, 16'd21323}; // indx = 3709
    #10;
    addra = 32'd118720;
    dina = {96'd0, 16'd3942, 16'd45978, 16'd56894, 16'd22667, 16'd57961, 16'd45178, 16'd58337, 16'd60280, 16'd31316, 16'd29341}; // indx = 3710
    #10;
    addra = 32'd118752;
    dina = {96'd0, 16'd32764, 16'd6658, 16'd22798, 16'd45215, 16'd36753, 16'd25929, 16'd31319, 16'd7514, 16'd18934, 16'd16421}; // indx = 3711
    #10;
    addra = 32'd118784;
    dina = {96'd0, 16'd54846, 16'd57320, 16'd41412, 16'd63925, 16'd10182, 16'd11626, 16'd26455, 16'd38009, 16'd58901, 16'd24033}; // indx = 3712
    #10;
    addra = 32'd118816;
    dina = {96'd0, 16'd11739, 16'd41150, 16'd45472, 16'd34148, 16'd43988, 16'd6241, 16'd20622, 16'd18535, 16'd36409, 16'd52334}; // indx = 3713
    #10;
    addra = 32'd118848;
    dina = {96'd0, 16'd19484, 16'd56767, 16'd10553, 16'd15784, 16'd8032, 16'd45264, 16'd62866, 16'd59761, 16'd25227, 16'd28371}; // indx = 3714
    #10;
    addra = 32'd118880;
    dina = {96'd0, 16'd56568, 16'd47701, 16'd61180, 16'd30416, 16'd14116, 16'd58005, 16'd25487, 16'd34935, 16'd56857, 16'd29953}; // indx = 3715
    #10;
    addra = 32'd118912;
    dina = {96'd0, 16'd21643, 16'd49060, 16'd29256, 16'd49892, 16'd60490, 16'd46724, 16'd19260, 16'd19007, 16'd16344, 16'd53679}; // indx = 3716
    #10;
    addra = 32'd118944;
    dina = {96'd0, 16'd25984, 16'd10105, 16'd15156, 16'd127, 16'd1819, 16'd8955, 16'd6106, 16'd24443, 16'd8821, 16'd15065}; // indx = 3717
    #10;
    addra = 32'd118976;
    dina = {96'd0, 16'd10599, 16'd24831, 16'd27669, 16'd59944, 16'd14080, 16'd17979, 16'd8539, 16'd21445, 16'd43559, 16'd52298}; // indx = 3718
    #10;
    addra = 32'd119008;
    dina = {96'd0, 16'd4075, 16'd6172, 16'd35558, 16'd709, 16'd43476, 16'd1560, 16'd58005, 16'd25084, 16'd46690, 16'd7611}; // indx = 3719
    #10;
    addra = 32'd119040;
    dina = {96'd0, 16'd53220, 16'd10103, 16'd40548, 16'd34593, 16'd10599, 16'd34165, 16'd44666, 16'd2576, 16'd44861, 16'd7828}; // indx = 3720
    #10;
    addra = 32'd119072;
    dina = {96'd0, 16'd40494, 16'd57536, 16'd22520, 16'd15494, 16'd43414, 16'd26019, 16'd39500, 16'd33070, 16'd24502, 16'd15620}; // indx = 3721
    #10;
    addra = 32'd119104;
    dina = {96'd0, 16'd58734, 16'd25015, 16'd31360, 16'd52614, 16'd26170, 16'd6620, 16'd42916, 16'd20971, 16'd49177, 16'd38547}; // indx = 3722
    #10;
    addra = 32'd119136;
    dina = {96'd0, 16'd46880, 16'd58440, 16'd27223, 16'd42345, 16'd23781, 16'd19493, 16'd52532, 16'd4062, 16'd17096, 16'd58500}; // indx = 3723
    #10;
    addra = 32'd119168;
    dina = {96'd0, 16'd10738, 16'd15269, 16'd13592, 16'd48871, 16'd10976, 16'd7558, 16'd27642, 16'd46698, 16'd47782, 16'd10740}; // indx = 3724
    #10;
    addra = 32'd119200;
    dina = {96'd0, 16'd38511, 16'd44578, 16'd3645, 16'd24103, 16'd26943, 16'd13257, 16'd37836, 16'd29559, 16'd8613, 16'd18194}; // indx = 3725
    #10;
    addra = 32'd119232;
    dina = {96'd0, 16'd8261, 16'd40742, 16'd2727, 16'd8509, 16'd37232, 16'd64726, 16'd34878, 16'd65037, 16'd7729, 16'd60902}; // indx = 3726
    #10;
    addra = 32'd119264;
    dina = {96'd0, 16'd40654, 16'd49846, 16'd2481, 16'd26629, 16'd14230, 16'd56838, 16'd40970, 16'd36968, 16'd49509, 16'd51641}; // indx = 3727
    #10;
    addra = 32'd119296;
    dina = {96'd0, 16'd30551, 16'd58649, 16'd44285, 16'd53069, 16'd38503, 16'd28716, 16'd58723, 16'd43407, 16'd38933, 16'd59017}; // indx = 3728
    #10;
    addra = 32'd119328;
    dina = {96'd0, 16'd7211, 16'd19957, 16'd7341, 16'd18652, 16'd15847, 16'd26743, 16'd24326, 16'd42626, 16'd15848, 16'd39250}; // indx = 3729
    #10;
    addra = 32'd119360;
    dina = {96'd0, 16'd34219, 16'd28527, 16'd1051, 16'd16862, 16'd50244, 16'd38689, 16'd22236, 16'd54608, 16'd48753, 16'd23788}; // indx = 3730
    #10;
    addra = 32'd119392;
    dina = {96'd0, 16'd22002, 16'd31249, 16'd64322, 16'd31216, 16'd17977, 16'd40222, 16'd29915, 16'd12280, 16'd20023, 16'd112}; // indx = 3731
    #10;
    addra = 32'd119424;
    dina = {96'd0, 16'd30936, 16'd30755, 16'd32918, 16'd19690, 16'd45009, 16'd34291, 16'd27397, 16'd62913, 16'd57022, 16'd55828}; // indx = 3732
    #10;
    addra = 32'd119456;
    dina = {96'd0, 16'd54551, 16'd30953, 16'd27448, 16'd21736, 16'd62500, 16'd8409, 16'd9690, 16'd17794, 16'd6858, 16'd35699}; // indx = 3733
    #10;
    addra = 32'd119488;
    dina = {96'd0, 16'd47996, 16'd65335, 16'd30545, 16'd59579, 16'd43564, 16'd26226, 16'd38469, 16'd39199, 16'd22367, 16'd40720}; // indx = 3734
    #10;
    addra = 32'd119520;
    dina = {96'd0, 16'd29302, 16'd8869, 16'd28337, 16'd43703, 16'd43794, 16'd64923, 16'd30509, 16'd62144, 16'd23564, 16'd35844}; // indx = 3735
    #10;
    addra = 32'd119552;
    dina = {96'd0, 16'd317, 16'd15209, 16'd62545, 16'd54594, 16'd47358, 16'd22865, 16'd21410, 16'd4440, 16'd11211, 16'd60342}; // indx = 3736
    #10;
    addra = 32'd119584;
    dina = {96'd0, 16'd41999, 16'd36078, 16'd49550, 16'd26023, 16'd17688, 16'd6696, 16'd36493, 16'd22641, 16'd25519, 16'd45694}; // indx = 3737
    #10;
    addra = 32'd119616;
    dina = {96'd0, 16'd59, 16'd12049, 16'd48257, 16'd17975, 16'd29417, 16'd55969, 16'd44630, 16'd12817, 16'd23948, 16'd37747}; // indx = 3738
    #10;
    addra = 32'd119648;
    dina = {96'd0, 16'd59250, 16'd28467, 16'd11823, 16'd22584, 16'd40300, 16'd40548, 16'd64543, 16'd15078, 16'd14774, 16'd26660}; // indx = 3739
    #10;
    addra = 32'd119680;
    dina = {96'd0, 16'd37753, 16'd50262, 16'd20553, 16'd3532, 16'd17889, 16'd12913, 16'd64490, 16'd44582, 16'd17328, 16'd62125}; // indx = 3740
    #10;
    addra = 32'd119712;
    dina = {96'd0, 16'd53729, 16'd1993, 16'd3246, 16'd39788, 16'd56640, 16'd60756, 16'd44236, 16'd2810, 16'd19727, 16'd45449}; // indx = 3741
    #10;
    addra = 32'd119744;
    dina = {96'd0, 16'd58778, 16'd5662, 16'd42794, 16'd35739, 16'd19221, 16'd5457, 16'd33758, 16'd53641, 16'd15450, 16'd11423}; // indx = 3742
    #10;
    addra = 32'd119776;
    dina = {96'd0, 16'd44781, 16'd6988, 16'd54763, 16'd62109, 16'd30052, 16'd45318, 16'd7823, 16'd47248, 16'd33711, 16'd65391}; // indx = 3743
    #10;
    addra = 32'd119808;
    dina = {96'd0, 16'd14118, 16'd33711, 16'd38012, 16'd4659, 16'd43099, 16'd54400, 16'd54009, 16'd31002, 16'd62302, 16'd21961}; // indx = 3744
    #10;
    addra = 32'd119840;
    dina = {96'd0, 16'd34074, 16'd50056, 16'd1605, 16'd25877, 16'd11702, 16'd54195, 16'd25398, 16'd55890, 16'd14864, 16'd19020}; // indx = 3745
    #10;
    addra = 32'd119872;
    dina = {96'd0, 16'd19787, 16'd5715, 16'd25824, 16'd12187, 16'd50493, 16'd59743, 16'd37395, 16'd12174, 16'd18770, 16'd54253}; // indx = 3746
    #10;
    addra = 32'd119904;
    dina = {96'd0, 16'd12690, 16'd12521, 16'd24984, 16'd54908, 16'd16314, 16'd12838, 16'd27073, 16'd64504, 16'd26961, 16'd9238}; // indx = 3747
    #10;
    addra = 32'd119936;
    dina = {96'd0, 16'd6648, 16'd23119, 16'd19099, 16'd8770, 16'd30730, 16'd41898, 16'd53598, 16'd26834, 16'd27624, 16'd15335}; // indx = 3748
    #10;
    addra = 32'd119968;
    dina = {96'd0, 16'd3063, 16'd30661, 16'd62925, 16'd36599, 16'd6908, 16'd55302, 16'd51493, 16'd16728, 16'd7208, 16'd63635}; // indx = 3749
    #10;
    addra = 32'd120000;
    dina = {96'd0, 16'd22566, 16'd54983, 16'd43656, 16'd3714, 16'd48259, 16'd16041, 16'd25197, 16'd28802, 16'd36800, 16'd53530}; // indx = 3750
    #10;
    addra = 32'd120032;
    dina = {96'd0, 16'd42589, 16'd47023, 16'd63778, 16'd35503, 16'd19776, 16'd36724, 16'd56832, 16'd36785, 16'd41001, 16'd297}; // indx = 3751
    #10;
    addra = 32'd120064;
    dina = {96'd0, 16'd2295, 16'd21874, 16'd27675, 16'd62595, 16'd43839, 16'd6442, 16'd10900, 16'd58462, 16'd909, 16'd53785}; // indx = 3752
    #10;
    addra = 32'd120096;
    dina = {96'd0, 16'd6461, 16'd36424, 16'd115, 16'd18541, 16'd5555, 16'd61354, 16'd20400, 16'd54162, 16'd13689, 16'd58554}; // indx = 3753
    #10;
    addra = 32'd120128;
    dina = {96'd0, 16'd17454, 16'd9612, 16'd3501, 16'd3003, 16'd47649, 16'd3594, 16'd32722, 16'd24493, 16'd13154, 16'd13582}; // indx = 3754
    #10;
    addra = 32'd120160;
    dina = {96'd0, 16'd23508, 16'd26638, 16'd43800, 16'd32817, 16'd64541, 16'd42594, 16'd32428, 16'd53478, 16'd9944, 16'd47050}; // indx = 3755
    #10;
    addra = 32'd120192;
    dina = {96'd0, 16'd36393, 16'd37245, 16'd10052, 16'd64376, 16'd22916, 16'd37814, 16'd21102, 16'd2141, 16'd41576, 16'd25489}; // indx = 3756
    #10;
    addra = 32'd120224;
    dina = {96'd0, 16'd40352, 16'd60160, 16'd21676, 16'd63561, 16'd13668, 16'd10283, 16'd3011, 16'd46016, 16'd37, 16'd40589}; // indx = 3757
    #10;
    addra = 32'd120256;
    dina = {96'd0, 16'd16492, 16'd7442, 16'd53723, 16'd31648, 16'd50072, 16'd19262, 16'd33185, 16'd9593, 16'd5434, 16'd29844}; // indx = 3758
    #10;
    addra = 32'd120288;
    dina = {96'd0, 16'd42502, 16'd41256, 16'd4368, 16'd52936, 16'd49769, 16'd13497, 16'd37833, 16'd28690, 16'd26838, 16'd30032}; // indx = 3759
    #10;
    addra = 32'd120320;
    dina = {96'd0, 16'd59691, 16'd31483, 16'd61100, 16'd54161, 16'd45264, 16'd20771, 16'd61460, 16'd42481, 16'd52792, 16'd31596}; // indx = 3760
    #10;
    addra = 32'd120352;
    dina = {96'd0, 16'd21961, 16'd61493, 16'd32939, 16'd29404, 16'd5178, 16'd57976, 16'd65027, 16'd9544, 16'd62241, 16'd41054}; // indx = 3761
    #10;
    addra = 32'd120384;
    dina = {96'd0, 16'd37488, 16'd27784, 16'd9324, 16'd21024, 16'd60793, 16'd16441, 16'd44733, 16'd933, 16'd7624, 16'd18086}; // indx = 3762
    #10;
    addra = 32'd120416;
    dina = {96'd0, 16'd16896, 16'd11422, 16'd36624, 16'd42289, 16'd29366, 16'd11200, 16'd43577, 16'd62944, 16'd5193, 16'd12505}; // indx = 3763
    #10;
    addra = 32'd120448;
    dina = {96'd0, 16'd64618, 16'd1345, 16'd3117, 16'd57522, 16'd45605, 16'd1053, 16'd19396, 16'd31070, 16'd7722, 16'd41301}; // indx = 3764
    #10;
    addra = 32'd120480;
    dina = {96'd0, 16'd16969, 16'd1116, 16'd9713, 16'd44098, 16'd42085, 16'd24092, 16'd29025, 16'd22340, 16'd41005, 16'd30473}; // indx = 3765
    #10;
    addra = 32'd120512;
    dina = {96'd0, 16'd22346, 16'd17259, 16'd19683, 16'd29084, 16'd3331, 16'd47681, 16'd23053, 16'd37904, 16'd39422, 16'd46988}; // indx = 3766
    #10;
    addra = 32'd120544;
    dina = {96'd0, 16'd24767, 16'd51069, 16'd60624, 16'd8972, 16'd41492, 16'd33414, 16'd28753, 16'd22263, 16'd20171, 16'd8851}; // indx = 3767
    #10;
    addra = 32'd120576;
    dina = {96'd0, 16'd15757, 16'd29666, 16'd55398, 16'd61550, 16'd1227, 16'd48078, 16'd20054, 16'd47955, 16'd1524, 16'd2107}; // indx = 3768
    #10;
    addra = 32'd120608;
    dina = {96'd0, 16'd25412, 16'd59610, 16'd14354, 16'd55305, 16'd22247, 16'd54636, 16'd13097, 16'd37499, 16'd23931, 16'd6187}; // indx = 3769
    #10;
    addra = 32'd120640;
    dina = {96'd0, 16'd45013, 16'd12526, 16'd23870, 16'd1270, 16'd63457, 16'd56627, 16'd14586, 16'd16441, 16'd32603, 16'd24031}; // indx = 3770
    #10;
    addra = 32'd120672;
    dina = {96'd0, 16'd18495, 16'd46069, 16'd42012, 16'd5220, 16'd918, 16'd62242, 16'd6464, 16'd17511, 16'd52750, 16'd9910}; // indx = 3771
    #10;
    addra = 32'd120704;
    dina = {96'd0, 16'd24255, 16'd46531, 16'd51874, 16'd46125, 16'd40665, 16'd25220, 16'd44520, 16'd22205, 16'd38041, 16'd34542}; // indx = 3772
    #10;
    addra = 32'd120736;
    dina = {96'd0, 16'd43404, 16'd11646, 16'd28735, 16'd48943, 16'd14266, 16'd47848, 16'd5271, 16'd18148, 16'd18578, 16'd47937}; // indx = 3773
    #10;
    addra = 32'd120768;
    dina = {96'd0, 16'd38953, 16'd65427, 16'd32757, 16'd56222, 16'd55725, 16'd30334, 16'd54090, 16'd17470, 16'd14951, 16'd1700}; // indx = 3774
    #10;
    addra = 32'd120800;
    dina = {96'd0, 16'd50868, 16'd23768, 16'd29726, 16'd28138, 16'd48033, 16'd56772, 16'd22546, 16'd49033, 16'd36494, 16'd45858}; // indx = 3775
    #10;
    addra = 32'd120832;
    dina = {96'd0, 16'd29662, 16'd56351, 16'd26375, 16'd22265, 16'd57192, 16'd3535, 16'd29481, 16'd59821, 16'd1721, 16'd2344}; // indx = 3776
    #10;
    addra = 32'd120864;
    dina = {96'd0, 16'd51893, 16'd54804, 16'd48007, 16'd20076, 16'd11511, 16'd2668, 16'd63175, 16'd45195, 16'd43914, 16'd34867}; // indx = 3777
    #10;
    addra = 32'd120896;
    dina = {96'd0, 16'd39861, 16'd38811, 16'd26731, 16'd5770, 16'd62417, 16'd64599, 16'd9762, 16'd2722, 16'd17888, 16'd53982}; // indx = 3778
    #10;
    addra = 32'd120928;
    dina = {96'd0, 16'd49856, 16'd40046, 16'd5537, 16'd62479, 16'd38499, 16'd30879, 16'd7018, 16'd26190, 16'd50561, 16'd11504}; // indx = 3779
    #10;
    addra = 32'd120960;
    dina = {96'd0, 16'd2663, 16'd779, 16'd33967, 16'd4256, 16'd10300, 16'd64867, 16'd46835, 16'd29607, 16'd51275, 16'd22458}; // indx = 3780
    #10;
    addra = 32'd120992;
    dina = {96'd0, 16'd51003, 16'd20996, 16'd43420, 16'd33403, 16'd4090, 16'd10535, 16'd42013, 16'd30049, 16'd49800, 16'd39687}; // indx = 3781
    #10;
    addra = 32'd121024;
    dina = {96'd0, 16'd34057, 16'd761, 16'd57519, 16'd54220, 16'd36152, 16'd56596, 16'd57360, 16'd13672, 16'd29689, 16'd50667}; // indx = 3782
    #10;
    addra = 32'd121056;
    dina = {96'd0, 16'd21497, 16'd26888, 16'd14194, 16'd18369, 16'd29273, 16'd52661, 16'd56088, 16'd48004, 16'd39853, 16'd23914}; // indx = 3783
    #10;
    addra = 32'd121088;
    dina = {96'd0, 16'd2332, 16'd48354, 16'd30236, 16'd6295, 16'd25759, 16'd5951, 16'd50187, 16'd21185, 16'd38718, 16'd52976}; // indx = 3784
    #10;
    addra = 32'd121120;
    dina = {96'd0, 16'd37800, 16'd29953, 16'd8349, 16'd14057, 16'd15928, 16'd58094, 16'd59802, 16'd52033, 16'd8012, 16'd16087}; // indx = 3785
    #10;
    addra = 32'd121152;
    dina = {96'd0, 16'd16633, 16'd59111, 16'd51121, 16'd28794, 16'd42642, 16'd64334, 16'd4751, 16'd51998, 16'd65379, 16'd57954}; // indx = 3786
    #10;
    addra = 32'd121184;
    dina = {96'd0, 16'd17517, 16'd62886, 16'd24889, 16'd41858, 16'd17898, 16'd56354, 16'd35312, 16'd2700, 16'd49781, 16'd30401}; // indx = 3787
    #10;
    addra = 32'd121216;
    dina = {96'd0, 16'd9804, 16'd48653, 16'd8675, 16'd12467, 16'd46657, 16'd23665, 16'd13613, 16'd58421, 16'd40288, 16'd30180}; // indx = 3788
    #10;
    addra = 32'd121248;
    dina = {96'd0, 16'd48629, 16'd64972, 16'd23886, 16'd39720, 16'd55928, 16'd57304, 16'd11208, 16'd1746, 16'd29690, 16'd50999}; // indx = 3789
    #10;
    addra = 32'd121280;
    dina = {96'd0, 16'd33648, 16'd36635, 16'd26622, 16'd56118, 16'd47306, 16'd13545, 16'd22621, 16'd10583, 16'd25251, 16'd47735}; // indx = 3790
    #10;
    addra = 32'd121312;
    dina = {96'd0, 16'd23204, 16'd25326, 16'd57639, 16'd41630, 16'd45791, 16'd61738, 16'd51777, 16'd44547, 16'd53085, 16'd60217}; // indx = 3791
    #10;
    addra = 32'd121344;
    dina = {96'd0, 16'd61086, 16'd43044, 16'd61140, 16'd55564, 16'd40849, 16'd34485, 16'd43061, 16'd48403, 16'd61401, 16'd65300}; // indx = 3792
    #10;
    addra = 32'd121376;
    dina = {96'd0, 16'd50591, 16'd21566, 16'd40448, 16'd41426, 16'd59943, 16'd60803, 16'd20804, 16'd38280, 16'd28368, 16'd4303}; // indx = 3793
    #10;
    addra = 32'd121408;
    dina = {96'd0, 16'd32494, 16'd45240, 16'd1901, 16'd227, 16'd27941, 16'd42131, 16'd63288, 16'd48460, 16'd18533, 16'd20468}; // indx = 3794
    #10;
    addra = 32'd121440;
    dina = {96'd0, 16'd16722, 16'd9026, 16'd15203, 16'd56898, 16'd55, 16'd4737, 16'd28549, 16'd23852, 16'd40239, 16'd6440}; // indx = 3795
    #10;
    addra = 32'd121472;
    dina = {96'd0, 16'd46705, 16'd15456, 16'd16340, 16'd26688, 16'd14313, 16'd18441, 16'd15516, 16'd40729, 16'd42181, 16'd7230}; // indx = 3796
    #10;
    addra = 32'd121504;
    dina = {96'd0, 16'd29291, 16'd45774, 16'd30455, 16'd52416, 16'd52564, 16'd32285, 16'd42106, 16'd5463, 16'd61839, 16'd48400}; // indx = 3797
    #10;
    addra = 32'd121536;
    dina = {96'd0, 16'd5839, 16'd40768, 16'd54603, 16'd18106, 16'd27495, 16'd33385, 16'd19088, 16'd9273, 16'd37993, 16'd27407}; // indx = 3798
    #10;
    addra = 32'd121568;
    dina = {96'd0, 16'd51719, 16'd49063, 16'd60690, 16'd19057, 16'd36370, 16'd52514, 16'd51771, 16'd7810, 16'd31427, 16'd49428}; // indx = 3799
    #10;
    addra = 32'd121600;
    dina = {96'd0, 16'd37507, 16'd37962, 16'd18703, 16'd45609, 16'd14326, 16'd16778, 16'd36485, 16'd50947, 16'd21013, 16'd43494}; // indx = 3800
    #10;
    addra = 32'd121632;
    dina = {96'd0, 16'd53011, 16'd1317, 16'd39889, 16'd896, 16'd45410, 16'd64573, 16'd47205, 16'd16977, 16'd56699, 16'd20039}; // indx = 3801
    #10;
    addra = 32'd121664;
    dina = {96'd0, 16'd25386, 16'd44166, 16'd7857, 16'd9993, 16'd22453, 16'd61344, 16'd64150, 16'd50514, 16'd23895, 16'd44912}; // indx = 3802
    #10;
    addra = 32'd121696;
    dina = {96'd0, 16'd64011, 16'd34506, 16'd64051, 16'd43466, 16'd6782, 16'd54312, 16'd32406, 16'd31998, 16'd15663, 16'd1392}; // indx = 3803
    #10;
    addra = 32'd121728;
    dina = {96'd0, 16'd3880, 16'd43457, 16'd18038, 16'd36971, 16'd24501, 16'd36263, 16'd54209, 16'd23908, 16'd49761, 16'd7280}; // indx = 3804
    #10;
    addra = 32'd121760;
    dina = {96'd0, 16'd20630, 16'd28802, 16'd46221, 16'd41891, 16'd21295, 16'd11039, 16'd42500, 16'd34327, 16'd8999, 16'd7644}; // indx = 3805
    #10;
    addra = 32'd121792;
    dina = {96'd0, 16'd53482, 16'd27089, 16'd38149, 16'd38929, 16'd43158, 16'd37282, 16'd8008, 16'd16175, 16'd12645, 16'd36376}; // indx = 3806
    #10;
    addra = 32'd121824;
    dina = {96'd0, 16'd58331, 16'd47369, 16'd39430, 16'd13348, 16'd52727, 16'd1298, 16'd60218, 16'd46080, 16'd28316, 16'd17340}; // indx = 3807
    #10;
    addra = 32'd121856;
    dina = {96'd0, 16'd18507, 16'd7323, 16'd5459, 16'd29762, 16'd55558, 16'd54503, 16'd2689, 16'd279, 16'd42721, 16'd662}; // indx = 3808
    #10;
    addra = 32'd121888;
    dina = {96'd0, 16'd27370, 16'd44731, 16'd41509, 16'd41768, 16'd62905, 16'd6797, 16'd9346, 16'd49397, 16'd61845, 16'd51991}; // indx = 3809
    #10;
    addra = 32'd121920;
    dina = {96'd0, 16'd2487, 16'd11535, 16'd61923, 16'd44441, 16'd36705, 16'd55508, 16'd54577, 16'd4231, 16'd32350, 16'd45195}; // indx = 3810
    #10;
    addra = 32'd121952;
    dina = {96'd0, 16'd33528, 16'd47986, 16'd48403, 16'd18672, 16'd32892, 16'd47756, 16'd7967, 16'd30295, 16'd58576, 16'd29487}; // indx = 3811
    #10;
    addra = 32'd121984;
    dina = {96'd0, 16'd1309, 16'd5347, 16'd19606, 16'd55708, 16'd22006, 16'd14209, 16'd8495, 16'd61240, 16'd45330, 16'd19243}; // indx = 3812
    #10;
    addra = 32'd122016;
    dina = {96'd0, 16'd20015, 16'd24512, 16'd10752, 16'd63956, 16'd62725, 16'd40409, 16'd62944, 16'd17558, 16'd6241, 16'd27770}; // indx = 3813
    #10;
    addra = 32'd122048;
    dina = {96'd0, 16'd62048, 16'd57993, 16'd17923, 16'd24675, 16'd41122, 16'd42893, 16'd32912, 16'd55342, 16'd55097, 16'd33062}; // indx = 3814
    #10;
    addra = 32'd122080;
    dina = {96'd0, 16'd29158, 16'd28983, 16'd31437, 16'd47376, 16'd58817, 16'd30107, 16'd51111, 16'd12598, 16'd63136, 16'd56969}; // indx = 3815
    #10;
    addra = 32'd122112;
    dina = {96'd0, 16'd56294, 16'd27855, 16'd29992, 16'd44592, 16'd20945, 16'd49526, 16'd31302, 16'd28424, 16'd487, 16'd32894}; // indx = 3816
    #10;
    addra = 32'd122144;
    dina = {96'd0, 16'd15002, 16'd42895, 16'd41125, 16'd56, 16'd40453, 16'd60150, 16'd7291, 16'd33991, 16'd63225, 16'd49397}; // indx = 3817
    #10;
    addra = 32'd122176;
    dina = {96'd0, 16'd3117, 16'd63896, 16'd4213, 16'd4923, 16'd15854, 16'd41246, 16'd8294, 16'd20933, 16'd3494, 16'd12858}; // indx = 3818
    #10;
    addra = 32'd122208;
    dina = {96'd0, 16'd33407, 16'd58138, 16'd56715, 16'd24500, 16'd20145, 16'd12388, 16'd36073, 16'd2669, 16'd26583, 16'd56512}; // indx = 3819
    #10;
    addra = 32'd122240;
    dina = {96'd0, 16'd63918, 16'd64957, 16'd25035, 16'd33829, 16'd39514, 16'd30845, 16'd2991, 16'd18674, 16'd16206, 16'd17827}; // indx = 3820
    #10;
    addra = 32'd122272;
    dina = {96'd0, 16'd49456, 16'd61948, 16'd27879, 16'd61494, 16'd28656, 16'd29326, 16'd31848, 16'd32670, 16'd46986, 16'd32187}; // indx = 3821
    #10;
    addra = 32'd122304;
    dina = {96'd0, 16'd8897, 16'd29416, 16'd43174, 16'd31606, 16'd39925, 16'd38628, 16'd36995, 16'd52379, 16'd28153, 16'd5990}; // indx = 3822
    #10;
    addra = 32'd122336;
    dina = {96'd0, 16'd36038, 16'd15701, 16'd15513, 16'd22799, 16'd20447, 16'd51802, 16'd50259, 16'd6689, 16'd48795, 16'd25944}; // indx = 3823
    #10;
    addra = 32'd122368;
    dina = {96'd0, 16'd42119, 16'd5267, 16'd48094, 16'd60408, 16'd33642, 16'd44196, 16'd12215, 16'd11595, 16'd61822, 16'd61328}; // indx = 3824
    #10;
    addra = 32'd122400;
    dina = {96'd0, 16'd16071, 16'd20656, 16'd29745, 16'd57570, 16'd32170, 16'd53173, 16'd7061, 16'd41491, 16'd18406, 16'd48440}; // indx = 3825
    #10;
    addra = 32'd122432;
    dina = {96'd0, 16'd39760, 16'd19142, 16'd20910, 16'd34815, 16'd3630, 16'd59145, 16'd3144, 16'd16699, 16'd52143, 16'd37808}; // indx = 3826
    #10;
    addra = 32'd122464;
    dina = {96'd0, 16'd5304, 16'd16597, 16'd55684, 16'd33888, 16'd7105, 16'd38983, 16'd9911, 16'd2542, 16'd25959, 16'd51179}; // indx = 3827
    #10;
    addra = 32'd122496;
    dina = {96'd0, 16'd20586, 16'd6679, 16'd64280, 16'd56182, 16'd43447, 16'd54689, 16'd5687, 16'd5980, 16'd13787, 16'd44793}; // indx = 3828
    #10;
    addra = 32'd122528;
    dina = {96'd0, 16'd29078, 16'd64820, 16'd27299, 16'd62271, 16'd2444, 16'd46718, 16'd29882, 16'd16470, 16'd34848, 16'd3618}; // indx = 3829
    #10;
    addra = 32'd122560;
    dina = {96'd0, 16'd54544, 16'd52784, 16'd38368, 16'd33128, 16'd43224, 16'd40412, 16'd47785, 16'd2227, 16'd42574, 16'd7746}; // indx = 3830
    #10;
    addra = 32'd122592;
    dina = {96'd0, 16'd28516, 16'd26929, 16'd24029, 16'd3178, 16'd64354, 16'd54684, 16'd45792, 16'd61703, 16'd17160, 16'd65513}; // indx = 3831
    #10;
    addra = 32'd122624;
    dina = {96'd0, 16'd18231, 16'd31938, 16'd13436, 16'd43369, 16'd9160, 16'd52253, 16'd32100, 16'd58491, 16'd31698, 16'd36488}; // indx = 3832
    #10;
    addra = 32'd122656;
    dina = {96'd0, 16'd1567, 16'd10195, 16'd12775, 16'd63320, 16'd45176, 16'd4508, 16'd3283, 16'd14202, 16'd56435, 16'd59172}; // indx = 3833
    #10;
    addra = 32'd122688;
    dina = {96'd0, 16'd28594, 16'd33646, 16'd36994, 16'd12251, 16'd60810, 16'd53751, 16'd39836, 16'd9000, 16'd61498, 16'd5273}; // indx = 3834
    #10;
    addra = 32'd122720;
    dina = {96'd0, 16'd22171, 16'd40856, 16'd2779, 16'd61639, 16'd15435, 16'd51763, 16'd10412, 16'd52396, 16'd2399, 16'd56442}; // indx = 3835
    #10;
    addra = 32'd122752;
    dina = {96'd0, 16'd47379, 16'd47143, 16'd63784, 16'd52589, 16'd13527, 16'd59491, 16'd8874, 16'd31997, 16'd49052, 16'd54406}; // indx = 3836
    #10;
    addra = 32'd122784;
    dina = {96'd0, 16'd25615, 16'd50641, 16'd29676, 16'd1142, 16'd24085, 16'd52355, 16'd8588, 16'd13152, 16'd15575, 16'd22626}; // indx = 3837
    #10;
    addra = 32'd122816;
    dina = {96'd0, 16'd61928, 16'd42077, 16'd840, 16'd56494, 16'd5624, 16'd45130, 16'd60723, 16'd56154, 16'd46619, 16'd20815}; // indx = 3838
    #10;
    addra = 32'd122848;
    dina = {96'd0, 16'd47513, 16'd14060, 16'd65530, 16'd10560, 16'd28856, 16'd33188, 16'd26114, 16'd53303, 16'd49496, 16'd58523}; // indx = 3839
    #10;
    addra = 32'd122880;
    dina = {96'd0, 16'd33212, 16'd35134, 16'd5026, 16'd10880, 16'd46317, 16'd19377, 16'd20607, 16'd36549, 16'd15969, 16'd53120}; // indx = 3840
    #10;
    addra = 32'd122912;
    dina = {96'd0, 16'd26305, 16'd10131, 16'd4783, 16'd50687, 16'd55820, 16'd20601, 16'd15966, 16'd31210, 16'd31413, 16'd30056}; // indx = 3841
    #10;
    addra = 32'd122944;
    dina = {96'd0, 16'd14129, 16'd45704, 16'd48428, 16'd7767, 16'd42968, 16'd34440, 16'd61463, 16'd9465, 16'd51069, 16'd33196}; // indx = 3842
    #10;
    addra = 32'd122976;
    dina = {96'd0, 16'd57610, 16'd36030, 16'd32659, 16'd19947, 16'd54208, 16'd30501, 16'd25274, 16'd40477, 16'd11913, 16'd16088}; // indx = 3843
    #10;
    addra = 32'd123008;
    dina = {96'd0, 16'd5935, 16'd34782, 16'd3552, 16'd13513, 16'd42488, 16'd16962, 16'd2762, 16'd29006, 16'd57691, 16'd23585}; // indx = 3844
    #10;
    addra = 32'd123040;
    dina = {96'd0, 16'd2958, 16'd14083, 16'd20182, 16'd51480, 16'd19076, 16'd62844, 16'd18133, 16'd13535, 16'd8425, 16'd54407}; // indx = 3845
    #10;
    addra = 32'd123072;
    dina = {96'd0, 16'd52754, 16'd3255, 16'd15679, 16'd50147, 16'd54173, 16'd13902, 16'd62831, 16'd26774, 16'd8277, 16'd62341}; // indx = 3846
    #10;
    addra = 32'd123104;
    dina = {96'd0, 16'd47302, 16'd2089, 16'd59448, 16'd645, 16'd36076, 16'd39989, 16'd28330, 16'd63073, 16'd30028, 16'd58992}; // indx = 3847
    #10;
    addra = 32'd123136;
    dina = {96'd0, 16'd41880, 16'd843, 16'd35267, 16'd10369, 16'd55891, 16'd14495, 16'd64864, 16'd35745, 16'd2442, 16'd44543}; // indx = 3848
    #10;
    addra = 32'd123168;
    dina = {96'd0, 16'd56258, 16'd11894, 16'd65438, 16'd10911, 16'd9134, 16'd31998, 16'd65509, 16'd21, 16'd9144, 16'd1951}; // indx = 3849
    #10;
    addra = 32'd123200;
    dina = {96'd0, 16'd32771, 16'd19886, 16'd16430, 16'd62507, 16'd13359, 16'd2917, 16'd32007, 16'd47290, 16'd60711, 16'd54674}; // indx = 3850
    #10;
    addra = 32'd123232;
    dina = {96'd0, 16'd36381, 16'd32934, 16'd13954, 16'd33294, 16'd40537, 16'd30036, 16'd59448, 16'd48804, 16'd64522, 16'd27411}; // indx = 3851
    #10;
    addra = 32'd123264;
    dina = {96'd0, 16'd16378, 16'd22646, 16'd3650, 16'd26544, 16'd60598, 16'd29839, 16'd2073, 16'd29869, 16'd61973, 16'd56364}; // indx = 3852
    #10;
    addra = 32'd123296;
    dina = {96'd0, 16'd28659, 16'd38429, 16'd24126, 16'd44071, 16'd58216, 16'd82, 16'd12726, 16'd63781, 16'd10387, 16'd31051}; // indx = 3853
    #10;
    addra = 32'd123328;
    dina = {96'd0, 16'd23003, 16'd29178, 16'd45998, 16'd11844, 16'd58012, 16'd24762, 16'd41288, 16'd472, 16'd39978, 16'd30864}; // indx = 3854
    #10;
    addra = 32'd123360;
    dina = {96'd0, 16'd27106, 16'd11324, 16'd53719, 16'd4662, 16'd44424, 16'd51218, 16'd10523, 16'd60604, 16'd14563, 16'd59465}; // indx = 3855
    #10;
    addra = 32'd123392;
    dina = {96'd0, 16'd7658, 16'd44717, 16'd58966, 16'd15120, 16'd47561, 16'd40688, 16'd41568, 16'd23193, 16'd4205, 16'd618}; // indx = 3856
    #10;
    addra = 32'd123424;
    dina = {96'd0, 16'd17280, 16'd62351, 16'd2525, 16'd30229, 16'd38703, 16'd31696, 16'd7228, 16'd26009, 16'd61568, 16'd14211}; // indx = 3857
    #10;
    addra = 32'd123456;
    dina = {96'd0, 16'd5342, 16'd55232, 16'd56777, 16'd46819, 16'd64456, 16'd50633, 16'd363, 16'd22867, 16'd9437, 16'd25322}; // indx = 3858
    #10;
    addra = 32'd123488;
    dina = {96'd0, 16'd55789, 16'd62081, 16'd5871, 16'd11549, 16'd6270, 16'd27239, 16'd14452, 16'd12141, 16'd3944, 16'd41777}; // indx = 3859
    #10;
    addra = 32'd123520;
    dina = {96'd0, 16'd16179, 16'd11172, 16'd40459, 16'd49294, 16'd13837, 16'd34788, 16'd43884, 16'd51271, 16'd41291, 16'd38248}; // indx = 3860
    #10;
    addra = 32'd123552;
    dina = {96'd0, 16'd37777, 16'd50940, 16'd18452, 16'd25144, 16'd4212, 16'd16303, 16'd60754, 16'd48855, 16'd50211, 16'd53556}; // indx = 3861
    #10;
    addra = 32'd123584;
    dina = {96'd0, 16'd55306, 16'd24247, 16'd45329, 16'd25010, 16'd43953, 16'd6869, 16'd60701, 16'd60684, 16'd30619, 16'd18351}; // indx = 3862
    #10;
    addra = 32'd123616;
    dina = {96'd0, 16'd25801, 16'd26915, 16'd36535, 16'd4906, 16'd55305, 16'd330, 16'd38309, 16'd54132, 16'd50521, 16'd5344}; // indx = 3863
    #10;
    addra = 32'd123648;
    dina = {96'd0, 16'd55958, 16'd48116, 16'd16457, 16'd25897, 16'd40383, 16'd52796, 16'd10893, 16'd42804, 16'd51161, 16'd57720}; // indx = 3864
    #10;
    addra = 32'd123680;
    dina = {96'd0, 16'd54769, 16'd33716, 16'd6565, 16'd59368, 16'd37324, 16'd41295, 16'd32676, 16'd54931, 16'd43378, 16'd37398}; // indx = 3865
    #10;
    addra = 32'd123712;
    dina = {96'd0, 16'd42528, 16'd30440, 16'd40302, 16'd58493, 16'd41731, 16'd14614, 16'd52237, 16'd23782, 16'd32274, 16'd41446}; // indx = 3866
    #10;
    addra = 32'd123744;
    dina = {96'd0, 16'd5188, 16'd17052, 16'd2634, 16'd17490, 16'd49617, 16'd20068, 16'd37541, 16'd19089, 16'd21882, 16'd38830}; // indx = 3867
    #10;
    addra = 32'd123776;
    dina = {96'd0, 16'd12900, 16'd46552, 16'd14946, 16'd57367, 16'd808, 16'd50259, 16'd22103, 16'd26111, 16'd16595, 16'd48487}; // indx = 3868
    #10;
    addra = 32'd123808;
    dina = {96'd0, 16'd59289, 16'd36387, 16'd26655, 16'd56647, 16'd25378, 16'd28423, 16'd22407, 16'd52279, 16'd17968, 16'd30727}; // indx = 3869
    #10;
    addra = 32'd123840;
    dina = {96'd0, 16'd50429, 16'd55276, 16'd54121, 16'd28075, 16'd37023, 16'd25241, 16'd63550, 16'd6242, 16'd44315, 16'd42262}; // indx = 3870
    #10;
    addra = 32'd123872;
    dina = {96'd0, 16'd27658, 16'd45966, 16'd20712, 16'd48335, 16'd43663, 16'd24875, 16'd55540, 16'd49520, 16'd830, 16'd58056}; // indx = 3871
    #10;
    addra = 32'd123904;
    dina = {96'd0, 16'd53129, 16'd55689, 16'd59429, 16'd50053, 16'd57874, 16'd49228, 16'd55569, 16'd3761, 16'd30366, 16'd61599}; // indx = 3872
    #10;
    addra = 32'd123936;
    dina = {96'd0, 16'd46429, 16'd22401, 16'd46771, 16'd62428, 16'd52374, 16'd47720, 16'd4054, 16'd24016, 16'd65043, 16'd28157}; // indx = 3873
    #10;
    addra = 32'd123968;
    dina = {96'd0, 16'd22663, 16'd38491, 16'd12963, 16'd19282, 16'd38112, 16'd51243, 16'd32107, 16'd28582, 16'd55135, 16'd59923}; // indx = 3874
    #10;
    addra = 32'd124000;
    dina = {96'd0, 16'd1752, 16'd13584, 16'd22601, 16'd47159, 16'd8359, 16'd13367, 16'd26787, 16'd22527, 16'd18717, 16'd59140}; // indx = 3875
    #10;
    addra = 32'd124032;
    dina = {96'd0, 16'd4547, 16'd51533, 16'd35673, 16'd51249, 16'd16609, 16'd60933, 16'd53813, 16'd32588, 16'd38772, 16'd4728}; // indx = 3876
    #10;
    addra = 32'd124064;
    dina = {96'd0, 16'd28541, 16'd25690, 16'd54863, 16'd20606, 16'd28542, 16'd12214, 16'd20191, 16'd29585, 16'd51412, 16'd26199}; // indx = 3877
    #10;
    addra = 32'd124096;
    dina = {96'd0, 16'd35640, 16'd7485, 16'd35439, 16'd23838, 16'd15124, 16'd20464, 16'd29103, 16'd30227, 16'd57702, 16'd43466}; // indx = 3878
    #10;
    addra = 32'd124128;
    dina = {96'd0, 16'd54374, 16'd5877, 16'd14447, 16'd2704, 16'd6904, 16'd42982, 16'd62596, 16'd15095, 16'd53262, 16'd8238}; // indx = 3879
    #10;
    addra = 32'd124160;
    dina = {96'd0, 16'd22243, 16'd61313, 16'd56114, 16'd9213, 16'd35958, 16'd53232, 16'd28303, 16'd53009, 16'd28332, 16'd63039}; // indx = 3880
    #10;
    addra = 32'd124192;
    dina = {96'd0, 16'd5176, 16'd29363, 16'd24202, 16'd611, 16'd51608, 16'd59854, 16'd62517, 16'd35367, 16'd29640, 16'd55904}; // indx = 3881
    #10;
    addra = 32'd124224;
    dina = {96'd0, 16'd55572, 16'd51126, 16'd34482, 16'd32313, 16'd5269, 16'd697, 16'd13457, 16'd1742, 16'd38893, 16'd21099}; // indx = 3882
    #10;
    addra = 32'd124256;
    dina = {96'd0, 16'd20655, 16'd15055, 16'd46476, 16'd44581, 16'd56667, 16'd63059, 16'd14171, 16'd22839, 16'd35389, 16'd15962}; // indx = 3883
    #10;
    addra = 32'd124288;
    dina = {96'd0, 16'd58900, 16'd44060, 16'd31515, 16'd37858, 16'd34322, 16'd23880, 16'd29985, 16'd11130, 16'd31868, 16'd21996}; // indx = 3884
    #10;
    addra = 32'd124320;
    dina = {96'd0, 16'd52138, 16'd63241, 16'd10998, 16'd36478, 16'd10433, 16'd28598, 16'd54351, 16'd39247, 16'd35300, 16'd64806}; // indx = 3885
    #10;
    addra = 32'd124352;
    dina = {96'd0, 16'd51920, 16'd26212, 16'd49807, 16'd10365, 16'd35063, 16'd30726, 16'd23510, 16'd62189, 16'd16704, 16'd45155}; // indx = 3886
    #10;
    addra = 32'd124384;
    dina = {96'd0, 16'd37295, 16'd32740, 16'd4141, 16'd19372, 16'd32764, 16'd52573, 16'd3915, 16'd4422, 16'd33436, 16'd26345}; // indx = 3887
    #10;
    addra = 32'd124416;
    dina = {96'd0, 16'd10686, 16'd15984, 16'd26202, 16'd10041, 16'd16174, 16'd64210, 16'd10975, 16'd14158, 16'd5331, 16'd29715}; // indx = 3888
    #10;
    addra = 32'd124448;
    dina = {96'd0, 16'd29909, 16'd887, 16'd2991, 16'd2056, 16'd40183, 16'd4603, 16'd36267, 16'd49782, 16'd56459, 16'd51507}; // indx = 3889
    #10;
    addra = 32'd124480;
    dina = {96'd0, 16'd20051, 16'd30245, 16'd58076, 16'd50695, 16'd26533, 16'd4648, 16'd8782, 16'd12911, 16'd39268, 16'd4277}; // indx = 3890
    #10;
    addra = 32'd124512;
    dina = {96'd0, 16'd7977, 16'd51070, 16'd23451, 16'd4236, 16'd15286, 16'd22639, 16'd10058, 16'd58493, 16'd46011, 16'd4595}; // indx = 3891
    #10;
    addra = 32'd124544;
    dina = {96'd0, 16'd38926, 16'd30563, 16'd18960, 16'd6297, 16'd839, 16'd64, 16'd4534, 16'd5139, 16'd53555, 16'd2705}; // indx = 3892
    #10;
    addra = 32'd124576;
    dina = {96'd0, 16'd19233, 16'd53172, 16'd41265, 16'd11296, 16'd11461, 16'd45629, 16'd16334, 16'd23860, 16'd26673, 16'd11244}; // indx = 3893
    #10;
    addra = 32'd124608;
    dina = {96'd0, 16'd40790, 16'd2930, 16'd41727, 16'd39013, 16'd36639, 16'd55058, 16'd38319, 16'd49433, 16'd53938, 16'd50955}; // indx = 3894
    #10;
    addra = 32'd124640;
    dina = {96'd0, 16'd39863, 16'd12020, 16'd19972, 16'd45563, 16'd48358, 16'd16416, 16'd45368, 16'd12028, 16'd44857, 16'd41885}; // indx = 3895
    #10;
    addra = 32'd124672;
    dina = {96'd0, 16'd23290, 16'd34557, 16'd32293, 16'd53737, 16'd5995, 16'd59200, 16'd29163, 16'd35551, 16'd38145, 16'd38411}; // indx = 3896
    #10;
    addra = 32'd124704;
    dina = {96'd0, 16'd51308, 16'd28923, 16'd3978, 16'd49342, 16'd24177, 16'd29297, 16'd58990, 16'd28128, 16'd8623, 16'd27843}; // indx = 3897
    #10;
    addra = 32'd124736;
    dina = {96'd0, 16'd64587, 16'd53063, 16'd55632, 16'd22200, 16'd13488, 16'd28338, 16'd48955, 16'd26104, 16'd34195, 16'd47768}; // indx = 3898
    #10;
    addra = 32'd124768;
    dina = {96'd0, 16'd489, 16'd292, 16'd14309, 16'd45409, 16'd30132, 16'd24731, 16'd52360, 16'd29796, 16'd17483, 16'd4729}; // indx = 3899
    #10;
    addra = 32'd124800;
    dina = {96'd0, 16'd12906, 16'd59548, 16'd55590, 16'd24440, 16'd22614, 16'd56606, 16'd36641, 16'd10761, 16'd6466, 16'd38130}; // indx = 3900
    #10;
    addra = 32'd124832;
    dina = {96'd0, 16'd6857, 16'd42330, 16'd20151, 16'd6002, 16'd25487, 16'd19450, 16'd34957, 16'd61435, 16'd65490, 16'd16387}; // indx = 3901
    #10;
    addra = 32'd124864;
    dina = {96'd0, 16'd8208, 16'd3639, 16'd11325, 16'd39752, 16'd65316, 16'd54986, 16'd49296, 16'd23326, 16'd17684, 16'd32458}; // indx = 3902
    #10;
    addra = 32'd124896;
    dina = {96'd0, 16'd11334, 16'd3286, 16'd30446, 16'd62881, 16'd44913, 16'd35062, 16'd62157, 16'd28316, 16'd22622, 16'd61778}; // indx = 3903
    #10;
    addra = 32'd124928;
    dina = {96'd0, 16'd47685, 16'd23178, 16'd39700, 16'd13274, 16'd26870, 16'd44732, 16'd53768, 16'd60494, 16'd61807, 16'd24198}; // indx = 3904
    #10;
    addra = 32'd124960;
    dina = {96'd0, 16'd51537, 16'd5164, 16'd35482, 16'd10702, 16'd24594, 16'd16674, 16'd49455, 16'd63661, 16'd51253, 16'd26769}; // indx = 3905
    #10;
    addra = 32'd124992;
    dina = {96'd0, 16'd44592, 16'd56077, 16'd30104, 16'd31888, 16'd53041, 16'd32435, 16'd56823, 16'd37197, 16'd7146, 16'd47068}; // indx = 3906
    #10;
    addra = 32'd125024;
    dina = {96'd0, 16'd51923, 16'd52856, 16'd21800, 16'd43444, 16'd52135, 16'd23549, 16'd15287, 16'd17345, 16'd53661, 16'd26009}; // indx = 3907
    #10;
    addra = 32'd125056;
    dina = {96'd0, 16'd41825, 16'd54456, 16'd44482, 16'd2447, 16'd2518, 16'd23539, 16'd61323, 16'd6798, 16'd30841, 16'd18376}; // indx = 3908
    #10;
    addra = 32'd125088;
    dina = {96'd0, 16'd21481, 16'd29286, 16'd47345, 16'd53231, 16'd56076, 16'd46906, 16'd5677, 16'd29301, 16'd21218, 16'd61054}; // indx = 3909
    #10;
    addra = 32'd125120;
    dina = {96'd0, 16'd54717, 16'd52837, 16'd54602, 16'd36523, 16'd51606, 16'd4189, 16'd30903, 16'd25307, 16'd32117, 16'd20009}; // indx = 3910
    #10;
    addra = 32'd125152;
    dina = {96'd0, 16'd19713, 16'd18578, 16'd33445, 16'd63235, 16'd12030, 16'd45133, 16'd62057, 16'd7292, 16'd31949, 16'd21203}; // indx = 3911
    #10;
    addra = 32'd125184;
    dina = {96'd0, 16'd50907, 16'd30285, 16'd43314, 16'd457, 16'd36817, 16'd26421, 16'd12073, 16'd52059, 16'd57238, 16'd10506}; // indx = 3912
    #10;
    addra = 32'd125216;
    dina = {96'd0, 16'd22495, 16'd17023, 16'd12215, 16'd54459, 16'd25741, 16'd19545, 16'd55400, 16'd20292, 16'd19841, 16'd55850}; // indx = 3913
    #10;
    addra = 32'd125248;
    dina = {96'd0, 16'd24734, 16'd344, 16'd32681, 16'd11629, 16'd35116, 16'd8083, 16'd62369, 16'd12665, 16'd12171, 16'd56192}; // indx = 3914
    #10;
    addra = 32'd125280;
    dina = {96'd0, 16'd38867, 16'd35015, 16'd50997, 16'd57448, 16'd11930, 16'd12072, 16'd36421, 16'd53156, 16'd51222, 16'd15115}; // indx = 3915
    #10;
    addra = 32'd125312;
    dina = {96'd0, 16'd18200, 16'd30864, 16'd407, 16'd46522, 16'd10234, 16'd41665, 16'd45502, 16'd33415, 16'd51301, 16'd12883}; // indx = 3916
    #10;
    addra = 32'd125344;
    dina = {96'd0, 16'd3652, 16'd796, 16'd3127, 16'd35700, 16'd61045, 16'd44085, 16'd1945, 16'd65293, 16'd55188, 16'd24360}; // indx = 3917
    #10;
    addra = 32'd125376;
    dina = {96'd0, 16'd55613, 16'd21859, 16'd55802, 16'd24392, 16'd56538, 16'd28116, 16'd25905, 16'd28668, 16'd37496, 16'd55373}; // indx = 3918
    #10;
    addra = 32'd125408;
    dina = {96'd0, 16'd17145, 16'd1916, 16'd4675, 16'd46336, 16'd3338, 16'd45296, 16'd29569, 16'd60749, 16'd5351, 16'd48962}; // indx = 3919
    #10;
    addra = 32'd125440;
    dina = {96'd0, 16'd16544, 16'd51911, 16'd45382, 16'd28173, 16'd15763, 16'd28168, 16'd20635, 16'd54640, 16'd23563, 16'd30575}; // indx = 3920
    #10;
    addra = 32'd125472;
    dina = {96'd0, 16'd31995, 16'd59581, 16'd43918, 16'd58976, 16'd33808, 16'd40234, 16'd37020, 16'd11627, 16'd22536, 16'd40039}; // indx = 3921
    #10;
    addra = 32'd125504;
    dina = {96'd0, 16'd35893, 16'd48785, 16'd40376, 16'd32296, 16'd40194, 16'd10161, 16'd9586, 16'd3482, 16'd54980, 16'd28792}; // indx = 3922
    #10;
    addra = 32'd125536;
    dina = {96'd0, 16'd35271, 16'd29689, 16'd40200, 16'd38494, 16'd9367, 16'd56576, 16'd59288, 16'd30517, 16'd42198, 16'd5627}; // indx = 3923
    #10;
    addra = 32'd125568;
    dina = {96'd0, 16'd53239, 16'd22030, 16'd45137, 16'd21441, 16'd25503, 16'd8696, 16'd1407, 16'd31983, 16'd34936, 16'd36042}; // indx = 3924
    #10;
    addra = 32'd125600;
    dina = {96'd0, 16'd55583, 16'd7735, 16'd60466, 16'd55811, 16'd7535, 16'd15278, 16'd4844, 16'd7194, 16'd14206, 16'd8244}; // indx = 3925
    #10;
    addra = 32'd125632;
    dina = {96'd0, 16'd50719, 16'd17667, 16'd28125, 16'd22446, 16'd42897, 16'd13215, 16'd26685, 16'd6201, 16'd51415, 16'd64306}; // indx = 3926
    #10;
    addra = 32'd125664;
    dina = {96'd0, 16'd15630, 16'd45557, 16'd14544, 16'd656, 16'd49281, 16'd3042, 16'd18173, 16'd39196, 16'd38249, 16'd37010}; // indx = 3927
    #10;
    addra = 32'd125696;
    dina = {96'd0, 16'd22522, 16'd28654, 16'd8104, 16'd60723, 16'd45774, 16'd60744, 16'd45169, 16'd17968, 16'd1758, 16'd52018}; // indx = 3928
    #10;
    addra = 32'd125728;
    dina = {96'd0, 16'd25332, 16'd29244, 16'd19795, 16'd15505, 16'd50038, 16'd38315, 16'd64146, 16'd37324, 16'd28692, 16'd32771}; // indx = 3929
    #10;
    addra = 32'd125760;
    dina = {96'd0, 16'd45814, 16'd20713, 16'd35909, 16'd58773, 16'd19018, 16'd1083, 16'd11999, 16'd43673, 16'd60143, 16'd55676}; // indx = 3930
    #10;
    addra = 32'd125792;
    dina = {96'd0, 16'd43719, 16'd40093, 16'd19287, 16'd32144, 16'd21482, 16'd60347, 16'd21843, 16'd27340, 16'd19626, 16'd49596}; // indx = 3931
    #10;
    addra = 32'd125824;
    dina = {96'd0, 16'd29480, 16'd54401, 16'd61926, 16'd9102, 16'd31819, 16'd28938, 16'd8673, 16'd22219, 16'd33303, 16'd44414}; // indx = 3932
    #10;
    addra = 32'd125856;
    dina = {96'd0, 16'd5941, 16'd41507, 16'd38015, 16'd61385, 16'd48215, 16'd38965, 16'd60840, 16'd4781, 16'd32105, 16'd7487}; // indx = 3933
    #10;
    addra = 32'd125888;
    dina = {96'd0, 16'd32615, 16'd60716, 16'd3909, 16'd2988, 16'd7930, 16'd5091, 16'd14468, 16'd38062, 16'd63456, 16'd55677}; // indx = 3934
    #10;
    addra = 32'd125920;
    dina = {96'd0, 16'd15922, 16'd10225, 16'd13769, 16'd32858, 16'd35144, 16'd1121, 16'd41043, 16'd38076, 16'd35593, 16'd29676}; // indx = 3935
    #10;
    addra = 32'd125952;
    dina = {96'd0, 16'd62348, 16'd40849, 16'd49140, 16'd9760, 16'd16104, 16'd32961, 16'd40140, 16'd45542, 16'd36238, 16'd64063}; // indx = 3936
    #10;
    addra = 32'd125984;
    dina = {96'd0, 16'd52112, 16'd12993, 16'd14920, 16'd36983, 16'd17863, 16'd37363, 16'd10529, 16'd31206, 16'd61655, 16'd14501}; // indx = 3937
    #10;
    addra = 32'd126016;
    dina = {96'd0, 16'd37989, 16'd59639, 16'd813, 16'd63306, 16'd13777, 16'd31044, 16'd30454, 16'd42774, 16'd34197, 16'd12793}; // indx = 3938
    #10;
    addra = 32'd126048;
    dina = {96'd0, 16'd11926, 16'd6027, 16'd12515, 16'd57865, 16'd18561, 16'd41133, 16'd60142, 16'd45159, 16'd7096, 16'd53861}; // indx = 3939
    #10;
    addra = 32'd126080;
    dina = {96'd0, 16'd7970, 16'd13991, 16'd48713, 16'd49444, 16'd24681, 16'd56187, 16'd48405, 16'd37744, 16'd6485, 16'd54717}; // indx = 3940
    #10;
    addra = 32'd126112;
    dina = {96'd0, 16'd59173, 16'd41748, 16'd62436, 16'd33110, 16'd43681, 16'd9183, 16'd57129, 16'd12617, 16'd37093, 16'd41648}; // indx = 3941
    #10;
    addra = 32'd126144;
    dina = {96'd0, 16'd12590, 16'd9518, 16'd17184, 16'd22417, 16'd53629, 16'd8249, 16'd36749, 16'd41289, 16'd10817, 16'd23676}; // indx = 3942
    #10;
    addra = 32'd126176;
    dina = {96'd0, 16'd50254, 16'd38002, 16'd4875, 16'd64819, 16'd39951, 16'd27912, 16'd10515, 16'd7922, 16'd3969, 16'd16618}; // indx = 3943
    #10;
    addra = 32'd126208;
    dina = {96'd0, 16'd28583, 16'd58827, 16'd14767, 16'd7007, 16'd60231, 16'd58166, 16'd57398, 16'd30156, 16'd21019, 16'd43130}; // indx = 3944
    #10;
    addra = 32'd126240;
    dina = {96'd0, 16'd47771, 16'd49116, 16'd38769, 16'd30229, 16'd29945, 16'd24060, 16'd6327, 16'd34246, 16'd51151, 16'd3295}; // indx = 3945
    #10;
    addra = 32'd126272;
    dina = {96'd0, 16'd32276, 16'd44722, 16'd42553, 16'd34173, 16'd40690, 16'd15518, 16'd20389, 16'd14590, 16'd29296, 16'd11261}; // indx = 3946
    #10;
    addra = 32'd126304;
    dina = {96'd0, 16'd31510, 16'd54358, 16'd9247, 16'd54227, 16'd30790, 16'd49539, 16'd7124, 16'd25880, 16'd2092, 16'd63133}; // indx = 3947
    #10;
    addra = 32'd126336;
    dina = {96'd0, 16'd29499, 16'd57671, 16'd14846, 16'd16358, 16'd33961, 16'd47229, 16'd41524, 16'd22555, 16'd65535, 16'd6116}; // indx = 3948
    #10;
    addra = 32'd126368;
    dina = {96'd0, 16'd1966, 16'd22981, 16'd12174, 16'd27216, 16'd23923, 16'd50069, 16'd49144, 16'd19113, 16'd11382, 16'd17842}; // indx = 3949
    #10;
    addra = 32'd126400;
    dina = {96'd0, 16'd59753, 16'd40145, 16'd14394, 16'd38104, 16'd40080, 16'd64365, 16'd4076, 16'd10796, 16'd40970, 16'd22010}; // indx = 3950
    #10;
    addra = 32'd126432;
    dina = {96'd0, 16'd58824, 16'd63750, 16'd42557, 16'd22071, 16'd10491, 16'd8643, 16'd16166, 16'd57991, 16'd39067, 16'd1205}; // indx = 3951
    #10;
    addra = 32'd126464;
    dina = {96'd0, 16'd56696, 16'd28189, 16'd45825, 16'd27069, 16'd48157, 16'd39906, 16'd45259, 16'd26008, 16'd15757, 16'd57389}; // indx = 3952
    #10;
    addra = 32'd126496;
    dina = {96'd0, 16'd50707, 16'd15454, 16'd43752, 16'd39807, 16'd10218, 16'd51872, 16'd58023, 16'd55617, 16'd58497, 16'd6606}; // indx = 3953
    #10;
    addra = 32'd126528;
    dina = {96'd0, 16'd45887, 16'd53563, 16'd18912, 16'd8573, 16'd44982, 16'd46461, 16'd57520, 16'd8826, 16'd59949, 16'd50317}; // indx = 3954
    #10;
    addra = 32'd126560;
    dina = {96'd0, 16'd5308, 16'd7696, 16'd58020, 16'd59321, 16'd50041, 16'd63411, 16'd4134, 16'd23834, 16'd48079, 16'd6868}; // indx = 3955
    #10;
    addra = 32'd126592;
    dina = {96'd0, 16'd6522, 16'd52404, 16'd56335, 16'd36859, 16'd55229, 16'd34465, 16'd40978, 16'd20977, 16'd12860, 16'd17942}; // indx = 3956
    #10;
    addra = 32'd126624;
    dina = {96'd0, 16'd12668, 16'd40409, 16'd5964, 16'd17581, 16'd28175, 16'd24465, 16'd51497, 16'd39806, 16'd41069, 16'd49203}; // indx = 3957
    #10;
    addra = 32'd126656;
    dina = {96'd0, 16'd9890, 16'd41366, 16'd41013, 16'd45655, 16'd52010, 16'd60143, 16'd50762, 16'd31501, 16'd2389, 16'd10549}; // indx = 3958
    #10;
    addra = 32'd126688;
    dina = {96'd0, 16'd22514, 16'd19165, 16'd24893, 16'd2825, 16'd15330, 16'd13362, 16'd18781, 16'd29374, 16'd44551, 16'd42648}; // indx = 3959
    #10;
    addra = 32'd126720;
    dina = {96'd0, 16'd60578, 16'd36705, 16'd12174, 16'd60672, 16'd53791, 16'd61356, 16'd18353, 16'd29860, 16'd2799, 16'd38944}; // indx = 3960
    #10;
    addra = 32'd126752;
    dina = {96'd0, 16'd11828, 16'd30052, 16'd1326, 16'd46448, 16'd43693, 16'd14720, 16'd27860, 16'd55860, 16'd3603, 16'd7715}; // indx = 3961
    #10;
    addra = 32'd126784;
    dina = {96'd0, 16'd2972, 16'd51292, 16'd20321, 16'd44269, 16'd27836, 16'd37084, 16'd1570, 16'd11283, 16'd54560, 16'd42234}; // indx = 3962
    #10;
    addra = 32'd126816;
    dina = {96'd0, 16'd13224, 16'd16142, 16'd58462, 16'd16640, 16'd20123, 16'd10651, 16'd1079, 16'd19339, 16'd26637, 16'd63489}; // indx = 3963
    #10;
    addra = 32'd126848;
    dina = {96'd0, 16'd60817, 16'd15440, 16'd51050, 16'd38356, 16'd62863, 16'd28843, 16'd14850, 16'd33297, 16'd3369, 16'd22598}; // indx = 3964
    #10;
    addra = 32'd126880;
    dina = {96'd0, 16'd39754, 16'd40370, 16'd61192, 16'd50201, 16'd10437, 16'd62328, 16'd1078, 16'd60872, 16'd13276, 16'd24630}; // indx = 3965
    #10;
    addra = 32'd126912;
    dina = {96'd0, 16'd46343, 16'd38700, 16'd61105, 16'd18210, 16'd39499, 16'd28666, 16'd34179, 16'd50779, 16'd18192, 16'd33148}; // indx = 3966
    #10;
    addra = 32'd126944;
    dina = {96'd0, 16'd39474, 16'd46490, 16'd2330, 16'd56145, 16'd610, 16'd3492, 16'd56529, 16'd29922, 16'd32119, 16'd10879}; // indx = 3967
    #10;
    addra = 32'd126976;
    dina = {96'd0, 16'd54762, 16'd7031, 16'd24914, 16'd53240, 16'd16808, 16'd18939, 16'd12886, 16'd10790, 16'd63279, 16'd844}; // indx = 3968
    #10;
    addra = 32'd127008;
    dina = {96'd0, 16'd50088, 16'd8174, 16'd265, 16'd33816, 16'd29059, 16'd21636, 16'd50287, 16'd64541, 16'd57161, 16'd25900}; // indx = 3969
    #10;
    addra = 32'd127040;
    dina = {96'd0, 16'd40661, 16'd22607, 16'd57843, 16'd10831, 16'd57661, 16'd10362, 16'd25935, 16'd50427, 16'd34240, 16'd2037}; // indx = 3970
    #10;
    addra = 32'd127072;
    dina = {96'd0, 16'd55964, 16'd55870, 16'd6313, 16'd33842, 16'd15071, 16'd47203, 16'd35233, 16'd25069, 16'd63896, 16'd2480}; // indx = 3971
    #10;
    addra = 32'd127104;
    dina = {96'd0, 16'd56650, 16'd9067, 16'd9798, 16'd8713, 16'd64767, 16'd46300, 16'd22595, 16'd50736, 16'd62984, 16'd45186}; // indx = 3972
    #10;
    addra = 32'd127136;
    dina = {96'd0, 16'd15331, 16'd42336, 16'd7271, 16'd39761, 16'd60239, 16'd41858, 16'd41352, 16'd4976, 16'd62267, 16'd43309}; // indx = 3973
    #10;
    addra = 32'd127168;
    dina = {96'd0, 16'd44097, 16'd54900, 16'd29062, 16'd28823, 16'd5965, 16'd37653, 16'd9448, 16'd39062, 16'd64078, 16'd58601}; // indx = 3974
    #10;
    addra = 32'd127200;
    dina = {96'd0, 16'd52745, 16'd14052, 16'd17610, 16'd47073, 16'd15468, 16'd12707, 16'd62755, 16'd23574, 16'd15122, 16'd40320}; // indx = 3975
    #10;
    addra = 32'd127232;
    dina = {96'd0, 16'd4088, 16'd60710, 16'd59016, 16'd14786, 16'd7137, 16'd57832, 16'd14170, 16'd4471, 16'd43533, 16'd59525}; // indx = 3976
    #10;
    addra = 32'd127264;
    dina = {96'd0, 16'd9716, 16'd59245, 16'd63940, 16'd31837, 16'd54211, 16'd40858, 16'd37202, 16'd35671, 16'd27749, 16'd61315}; // indx = 3977
    #10;
    addra = 32'd127296;
    dina = {96'd0, 16'd34756, 16'd41856, 16'd65476, 16'd35604, 16'd36012, 16'd32549, 16'd45895, 16'd62847, 16'd50777, 16'd29131}; // indx = 3978
    #10;
    addra = 32'd127328;
    dina = {96'd0, 16'd59664, 16'd59617, 16'd2360, 16'd23505, 16'd30691, 16'd18467, 16'd64885, 16'd44699, 16'd2053, 16'd15604}; // indx = 3979
    #10;
    addra = 32'd127360;
    dina = {96'd0, 16'd38315, 16'd45291, 16'd28072, 16'd60199, 16'd37581, 16'd32284, 16'd24530, 16'd20557, 16'd17204, 16'd45375}; // indx = 3980
    #10;
    addra = 32'd127392;
    dina = {96'd0, 16'd37466, 16'd53570, 16'd62822, 16'd59861, 16'd36010, 16'd24499, 16'd49530, 16'd5612, 16'd64712, 16'd37904}; // indx = 3981
    #10;
    addra = 32'd127424;
    dina = {96'd0, 16'd27876, 16'd53990, 16'd51465, 16'd49264, 16'd35229, 16'd2978, 16'd54559, 16'd44739, 16'd28556, 16'd6586}; // indx = 3982
    #10;
    addra = 32'd127456;
    dina = {96'd0, 16'd23013, 16'd57613, 16'd35459, 16'd40932, 16'd27267, 16'd4624, 16'd36600, 16'd34199, 16'd33525, 16'd18801}; // indx = 3983
    #10;
    addra = 32'd127488;
    dina = {96'd0, 16'd53091, 16'd4698, 16'd35374, 16'd12636, 16'd59412, 16'd49729, 16'd27210, 16'd1702, 16'd585, 16'd63321}; // indx = 3984
    #10;
    addra = 32'd127520;
    dina = {96'd0, 16'd57528, 16'd61501, 16'd43129, 16'd43382, 16'd48843, 16'd10737, 16'd46367, 16'd61131, 16'd34189, 16'd40319}; // indx = 3985
    #10;
    addra = 32'd127552;
    dina = {96'd0, 16'd11792, 16'd42019, 16'd37716, 16'd19633, 16'd47860, 16'd55967, 16'd47276, 16'd40034, 16'd50914, 16'd37436}; // indx = 3986
    #10;
    addra = 32'd127584;
    dina = {96'd0, 16'd10991, 16'd15937, 16'd10917, 16'd62141, 16'd16155, 16'd46643, 16'd33206, 16'd17658, 16'd17499, 16'd15539}; // indx = 3987
    #10;
    addra = 32'd127616;
    dina = {96'd0, 16'd6165, 16'd27494, 16'd52687, 16'd23291, 16'd28126, 16'd56111, 16'd48926, 16'd48471, 16'd44383, 16'd13552}; // indx = 3988
    #10;
    addra = 32'd127648;
    dina = {96'd0, 16'd30353, 16'd13755, 16'd27391, 16'd30636, 16'd46965, 16'd34508, 16'd9866, 16'd47384, 16'd28676, 16'd225}; // indx = 3989
    #10;
    addra = 32'd127680;
    dina = {96'd0, 16'd30667, 16'd5487, 16'd65101, 16'd49076, 16'd58505, 16'd43797, 16'd29879, 16'd45821, 16'd40601, 16'd64219}; // indx = 3990
    #10;
    addra = 32'd127712;
    dina = {96'd0, 16'd13518, 16'd55844, 16'd2984, 16'd55617, 16'd8390, 16'd15171, 16'd52470, 16'd1571, 16'd45513, 16'd51035}; // indx = 3991
    #10;
    addra = 32'd127744;
    dina = {96'd0, 16'd18659, 16'd45573, 16'd60660, 16'd5635, 16'd43853, 16'd37665, 16'd51777, 16'd8583, 16'd34351, 16'd34875}; // indx = 3992
    #10;
    addra = 32'd127776;
    dina = {96'd0, 16'd22351, 16'd21263, 16'd22523, 16'd52213, 16'd21550, 16'd31517, 16'd41284, 16'd33093, 16'd44094, 16'd38264}; // indx = 3993
    #10;
    addra = 32'd127808;
    dina = {96'd0, 16'd53205, 16'd18272, 16'd59794, 16'd12341, 16'd26827, 16'd2935, 16'd52028, 16'd55184, 16'd12297, 16'd26676}; // indx = 3994
    #10;
    addra = 32'd127840;
    dina = {96'd0, 16'd20475, 16'd38704, 16'd11408, 16'd23909, 16'd37586, 16'd6457, 16'd15017, 16'd39462, 16'd13252, 16'd58631}; // indx = 3995
    #10;
    addra = 32'd127872;
    dina = {96'd0, 16'd48319, 16'd41607, 16'd51652, 16'd43828, 16'd8750, 16'd62056, 16'd63846, 16'd28370, 16'd44009, 16'd56149}; // indx = 3996
    #10;
    addra = 32'd127904;
    dina = {96'd0, 16'd45234, 16'd8240, 16'd44229, 16'd9005, 16'd20180, 16'd50756, 16'd64489, 16'd14048, 16'd56978, 16'd42715}; // indx = 3997
    #10;
    addra = 32'd127936;
    dina = {96'd0, 16'd41324, 16'd9073, 16'd42516, 16'd21851, 16'd26421, 16'd52697, 16'd60975, 16'd57004, 16'd18647, 16'd22142}; // indx = 3998
    #10;
    addra = 32'd127968;
    dina = {96'd0, 16'd37524, 16'd40818, 16'd27991, 16'd13569, 16'd28244, 16'd14985, 16'd29144, 16'd8848, 16'd12644, 16'd36612}; // indx = 3999
    #10;
    addra = 32'd128000;
    dina = {96'd0, 16'd11680, 16'd45397, 16'd50381, 16'd40689, 16'd60457, 16'd59428, 16'd64174, 16'd6496, 16'd65293, 16'd16158}; // indx = 4000
    #10;
    addra = 32'd128032;
    dina = {96'd0, 16'd24248, 16'd38375, 16'd28278, 16'd11008, 16'd46344, 16'd23240, 16'd7053, 16'd14128, 16'd15221, 16'd40544}; // indx = 4001
    #10;
    addra = 32'd128064;
    dina = {96'd0, 16'd36840, 16'd44898, 16'd49801, 16'd52272, 16'd60760, 16'd23907, 16'd5486, 16'd60675, 16'd44016, 16'd2083}; // indx = 4002
    #10;
    addra = 32'd128096;
    dina = {96'd0, 16'd46342, 16'd40199, 16'd6196, 16'd58723, 16'd39254, 16'd17592, 16'd50295, 16'd40949, 16'd160, 16'd63693}; // indx = 4003
    #10;
    addra = 32'd128128;
    dina = {96'd0, 16'd64624, 16'd3330, 16'd47010, 16'd32889, 16'd58415, 16'd9750, 16'd7524, 16'd18489, 16'd1719, 16'd50839}; // indx = 4004
    #10;
    addra = 32'd128160;
    dina = {96'd0, 16'd13627, 16'd58509, 16'd41698, 16'd41909, 16'd17551, 16'd42438, 16'd63430, 16'd63012, 16'd12557, 16'd35960}; // indx = 4005
    #10;
    addra = 32'd128192;
    dina = {96'd0, 16'd35075, 16'd46170, 16'd17609, 16'd58993, 16'd55271, 16'd16196, 16'd45490, 16'd44718, 16'd24148, 16'd3255}; // indx = 4006
    #10;
    addra = 32'd128224;
    dina = {96'd0, 16'd49067, 16'd57785, 16'd53591, 16'd5019, 16'd14925, 16'd39675, 16'd27828, 16'd22221, 16'd42349, 16'd51740}; // indx = 4007
    #10;
    addra = 32'd128256;
    dina = {96'd0, 16'd12031, 16'd23602, 16'd18324, 16'd43486, 16'd65492, 16'd7089, 16'd64442, 16'd43778, 16'd40749, 16'd23936}; // indx = 4008
    #10;
    addra = 32'd128288;
    dina = {96'd0, 16'd60551, 16'd35123, 16'd23241, 16'd13891, 16'd520, 16'd27082, 16'd25356, 16'd26700, 16'd54426, 16'd39357}; // indx = 4009
    #10;
    addra = 32'd128320;
    dina = {96'd0, 16'd35914, 16'd58368, 16'd21319, 16'd19715, 16'd31753, 16'd53694, 16'd39099, 16'd51903, 16'd38020, 16'd31244}; // indx = 4010
    #10;
    addra = 32'd128352;
    dina = {96'd0, 16'd48240, 16'd24546, 16'd62107, 16'd6359, 16'd62091, 16'd47289, 16'd64655, 16'd41831, 16'd53952, 16'd43564}; // indx = 4011
    #10;
    addra = 32'd128384;
    dina = {96'd0, 16'd9716, 16'd7934, 16'd18859, 16'd35197, 16'd57399, 16'd15156, 16'd55573, 16'd35258, 16'd34294, 16'd60462}; // indx = 4012
    #10;
    addra = 32'd128416;
    dina = {96'd0, 16'd34223, 16'd14178, 16'd52424, 16'd33390, 16'd28429, 16'd35000, 16'd13117, 16'd58381, 16'd35038, 16'd8326}; // indx = 4013
    #10;
    addra = 32'd128448;
    dina = {96'd0, 16'd63751, 16'd35248, 16'd49629, 16'd13736, 16'd38272, 16'd29624, 16'd44206, 16'd62990, 16'd20961, 16'd7493}; // indx = 4014
    #10;
    addra = 32'd128480;
    dina = {96'd0, 16'd65065, 16'd29560, 16'd19417, 16'd61542, 16'd49920, 16'd60564, 16'd36078, 16'd51796, 16'd54641, 16'd55975}; // indx = 4015
    #10;
    addra = 32'd128512;
    dina = {96'd0, 16'd48724, 16'd36902, 16'd63849, 16'd51401, 16'd21578, 16'd35356, 16'd7605, 16'd61191, 16'd13596, 16'd33304}; // indx = 4016
    #10;
    addra = 32'd128544;
    dina = {96'd0, 16'd14729, 16'd10200, 16'd36008, 16'd20388, 16'd47828, 16'd61576, 16'd35387, 16'd47113, 16'd48947, 16'd53773}; // indx = 4017
    #10;
    addra = 32'd128576;
    dina = {96'd0, 16'd48428, 16'd16479, 16'd53215, 16'd41729, 16'd42385, 16'd30290, 16'd18865, 16'd64872, 16'd22316, 16'd12215}; // indx = 4018
    #10;
    addra = 32'd128608;
    dina = {96'd0, 16'd58995, 16'd5674, 16'd45438, 16'd58177, 16'd55148, 16'd53346, 16'd34558, 16'd63191, 16'd45674, 16'd58411}; // indx = 4019
    #10;
    addra = 32'd128640;
    dina = {96'd0, 16'd62814, 16'd41318, 16'd30186, 16'd56873, 16'd63260, 16'd61713, 16'd45405, 16'd7059, 16'd25325, 16'd61124}; // indx = 4020
    #10;
    addra = 32'd128672;
    dina = {96'd0, 16'd18367, 16'd37895, 16'd32707, 16'd38999, 16'd10589, 16'd53809, 16'd47095, 16'd40532, 16'd20460, 16'd8982}; // indx = 4021
    #10;
    addra = 32'd128704;
    dina = {96'd0, 16'd18715, 16'd19224, 16'd6347, 16'd26159, 16'd1921, 16'd35116, 16'd58587, 16'd29809, 16'd1251, 16'd30199}; // indx = 4022
    #10;
    addra = 32'd128736;
    dina = {96'd0, 16'd36710, 16'd31394, 16'd42184, 16'd38562, 16'd34772, 16'd2097, 16'd10926, 16'd27636, 16'd63892, 16'd19691}; // indx = 4023
    #10;
    addra = 32'd128768;
    dina = {96'd0, 16'd50288, 16'd53348, 16'd55127, 16'd58762, 16'd55504, 16'd47266, 16'd25599, 16'd22477, 16'd1892, 16'd41730}; // indx = 4024
    #10;
    addra = 32'd128800;
    dina = {96'd0, 16'd60570, 16'd11313, 16'd63438, 16'd26127, 16'd19267, 16'd42402, 16'd3067, 16'd60553, 16'd41770, 16'd58427}; // indx = 4025
    #10;
    addra = 32'd128832;
    dina = {96'd0, 16'd25814, 16'd36725, 16'd61844, 16'd44353, 16'd3170, 16'd527, 16'd28110, 16'd23635, 16'd6292, 16'd54697}; // indx = 4026
    #10;
    addra = 32'd128864;
    dina = {96'd0, 16'd37587, 16'd44094, 16'd64825, 16'd57430, 16'd34061, 16'd819, 16'd41947, 16'd62511, 16'd64418, 16'd56275}; // indx = 4027
    #10;
    addra = 32'd128896;
    dina = {96'd0, 16'd676, 16'd26327, 16'd18039, 16'd16178, 16'd42394, 16'd57845, 16'd56609, 16'd54985, 16'd45895, 16'd43816}; // indx = 4028
    #10;
    addra = 32'd128928;
    dina = {96'd0, 16'd51877, 16'd29415, 16'd25341, 16'd54574, 16'd45625, 16'd37083, 16'd56985, 16'd65257, 16'd12934, 16'd56855}; // indx = 4029
    #10;
    addra = 32'd128960;
    dina = {96'd0, 16'd43508, 16'd58276, 16'd42834, 16'd23970, 16'd10580, 16'd19499, 16'd61892, 16'd53608, 16'd27539, 16'd50469}; // indx = 4030
    #10;
    addra = 32'd128992;
    dina = {96'd0, 16'd44114, 16'd29558, 16'd60787, 16'd20868, 16'd20859, 16'd42685, 16'd49645, 16'd45190, 16'd59167, 16'd10559}; // indx = 4031
    #10;
    addra = 32'd129024;
    dina = {96'd0, 16'd17538, 16'd51319, 16'd47061, 16'd3799, 16'd56157, 16'd29013, 16'd52007, 16'd30519, 16'd25253, 16'd12448}; // indx = 4032
    #10;
    addra = 32'd129056;
    dina = {96'd0, 16'd25148, 16'd31839, 16'd60042, 16'd45842, 16'd3949, 16'd60966, 16'd22567, 16'd61551, 16'd46473, 16'd64685}; // indx = 4033
    #10;
    addra = 32'd129088;
    dina = {96'd0, 16'd47172, 16'd3117, 16'd33489, 16'd26032, 16'd37374, 16'd40642, 16'd33716, 16'd56574, 16'd30723, 16'd9388}; // indx = 4034
    #10;
    addra = 32'd129120;
    dina = {96'd0, 16'd25524, 16'd37869, 16'd44838, 16'd59973, 16'd40957, 16'd63601, 16'd8049, 16'd63080, 16'd49108, 16'd57777}; // indx = 4035
    #10;
    addra = 32'd129152;
    dina = {96'd0, 16'd20286, 16'd4788, 16'd9654, 16'd11611, 16'd43306, 16'd36072, 16'd54905, 16'd64544, 16'd9037, 16'd29823}; // indx = 4036
    #10;
    addra = 32'd129184;
    dina = {96'd0, 16'd37413, 16'd2174, 16'd62330, 16'd18690, 16'd51858, 16'd38999, 16'd4228, 16'd10971, 16'd9383, 16'd43292}; // indx = 4037
    #10;
    addra = 32'd129216;
    dina = {96'd0, 16'd55646, 16'd8499, 16'd51637, 16'd48680, 16'd65041, 16'd35626, 16'd21775, 16'd39844, 16'd29277, 16'd6246}; // indx = 4038
    #10;
    addra = 32'd129248;
    dina = {96'd0, 16'd48647, 16'd16395, 16'd17628, 16'd10839, 16'd10454, 16'd14996, 16'd21625, 16'd60343, 16'd64800, 16'd4562}; // indx = 4039
    #10;
    addra = 32'd129280;
    dina = {96'd0, 16'd2826, 16'd3241, 16'd46642, 16'd14786, 16'd25511, 16'd34267, 16'd21872, 16'd27802, 16'd26694, 16'd49427}; // indx = 4040
    #10;
    addra = 32'd129312;
    dina = {96'd0, 16'd50889, 16'd55456, 16'd5227, 16'd34386, 16'd11753, 16'd61413, 16'd45757, 16'd62881, 16'd39237, 16'd44073}; // indx = 4041
    #10;
    addra = 32'd129344;
    dina = {96'd0, 16'd55111, 16'd62923, 16'd49786, 16'd10589, 16'd62632, 16'd27369, 16'd34340, 16'd15488, 16'd12796, 16'd21990}; // indx = 4042
    #10;
    addra = 32'd129376;
    dina = {96'd0, 16'd29153, 16'd5170, 16'd27187, 16'd64657, 16'd46557, 16'd58990, 16'd41916, 16'd42075, 16'd14362, 16'd54738}; // indx = 4043
    #10;
    addra = 32'd129408;
    dina = {96'd0, 16'd34337, 16'd14236, 16'd63179, 16'd62710, 16'd41679, 16'd30535, 16'd50946, 16'd9161, 16'd41266, 16'd25027}; // indx = 4044
    #10;
    addra = 32'd129440;
    dina = {96'd0, 16'd57128, 16'd3105, 16'd57397, 16'd10876, 16'd18144, 16'd37802, 16'd30404, 16'd41622, 16'd45930, 16'd28807}; // indx = 4045
    #10;
    addra = 32'd129472;
    dina = {96'd0, 16'd13395, 16'd13741, 16'd51224, 16'd47787, 16'd17165, 16'd47338, 16'd51277, 16'd21616, 16'd1547, 16'd51004}; // indx = 4046
    #10;
    addra = 32'd129504;
    dina = {96'd0, 16'd57525, 16'd44840, 16'd40280, 16'd33032, 16'd56297, 16'd51662, 16'd24487, 16'd7125, 16'd58274, 16'd44615}; // indx = 4047
    #10;
    addra = 32'd129536;
    dina = {96'd0, 16'd4025, 16'd26941, 16'd10777, 16'd14402, 16'd22291, 16'd60248, 16'd47538, 16'd56730, 16'd43627, 16'd20230}; // indx = 4048
    #10;
    addra = 32'd129568;
    dina = {96'd0, 16'd17401, 16'd32572, 16'd10822, 16'd26824, 16'd3462, 16'd19290, 16'd3419, 16'd44744, 16'd13012, 16'd14734}; // indx = 4049
    #10;
    addra = 32'd129600;
    dina = {96'd0, 16'd42257, 16'd31626, 16'd46764, 16'd27798, 16'd362, 16'd43825, 16'd61599, 16'd9464, 16'd49618, 16'd15217}; // indx = 4050
    #10;
    addra = 32'd129632;
    dina = {96'd0, 16'd63872, 16'd45465, 16'd19175, 16'd7670, 16'd56233, 16'd1874, 16'd60994, 16'd34441, 16'd58383, 16'd32809}; // indx = 4051
    #10;
    addra = 32'd129664;
    dina = {96'd0, 16'd48076, 16'd60952, 16'd36248, 16'd13321, 16'd50065, 16'd7934, 16'd16541, 16'd43402, 16'd48564, 16'd2538}; // indx = 4052
    #10;
    addra = 32'd129696;
    dina = {96'd0, 16'd380, 16'd9835, 16'd45238, 16'd56513, 16'd14070, 16'd8533, 16'd7111, 16'd17742, 16'd2642, 16'd4577}; // indx = 4053
    #10;
    addra = 32'd129728;
    dina = {96'd0, 16'd57365, 16'd23644, 16'd29265, 16'd21455, 16'd35792, 16'd17841, 16'd28902, 16'd39489, 16'd13029, 16'd55814}; // indx = 4054
    #10;
    addra = 32'd129760;
    dina = {96'd0, 16'd21122, 16'd19724, 16'd14806, 16'd15362, 16'd18446, 16'd19184, 16'd37882, 16'd26821, 16'd41489, 16'd28207}; // indx = 4055
    #10;
    addra = 32'd129792;
    dina = {96'd0, 16'd62446, 16'd41069, 16'd14540, 16'd24363, 16'd30023, 16'd48476, 16'd18273, 16'd50121, 16'd31807, 16'd22008}; // indx = 4056
    #10;
    addra = 32'd129824;
    dina = {96'd0, 16'd57230, 16'd30115, 16'd65083, 16'd22340, 16'd30600, 16'd13872, 16'd51973, 16'd6366, 16'd30513, 16'd60235}; // indx = 4057
    #10;
    addra = 32'd129856;
    dina = {96'd0, 16'd52829, 16'd34402, 16'd52967, 16'd39554, 16'd16924, 16'd35066, 16'd18638, 16'd28958, 16'd59524, 16'd64924}; // indx = 4058
    #10;
    addra = 32'd129888;
    dina = {96'd0, 16'd43874, 16'd26570, 16'd37567, 16'd7287, 16'd26885, 16'd34747, 16'd54536, 16'd64712, 16'd61737, 16'd62090}; // indx = 4059
    #10;
    addra = 32'd129920;
    dina = {96'd0, 16'd41057, 16'd60949, 16'd49465, 16'd43421, 16'd21553, 16'd5174, 16'd11155, 16'd12504, 16'd59792, 16'd21908}; // indx = 4060
    #10;
    addra = 32'd129952;
    dina = {96'd0, 16'd40194, 16'd8175, 16'd35738, 16'd39759, 16'd21748, 16'd31670, 16'd58783, 16'd297, 16'd18567, 16'd9879}; // indx = 4061
    #10;
    addra = 32'd129984;
    dina = {96'd0, 16'd59113, 16'd2766, 16'd25439, 16'd29428, 16'd25987, 16'd62332, 16'd9166, 16'd63845, 16'd20656, 16'd22460}; // indx = 4062
    #10;
    addra = 32'd130016;
    dina = {96'd0, 16'd43415, 16'd42602, 16'd45746, 16'd25057, 16'd20331, 16'd54645, 16'd32691, 16'd10968, 16'd45449, 16'd63258}; // indx = 4063
    #10;
    addra = 32'd130048;
    dina = {96'd0, 16'd37673, 16'd49208, 16'd53453, 16'd39740, 16'd59506, 16'd3768, 16'd25261, 16'd29870, 16'd16098, 16'd17125}; // indx = 4064
    #10;
    addra = 32'd130080;
    dina = {96'd0, 16'd5498, 16'd39641, 16'd9594, 16'd33719, 16'd65279, 16'd49423, 16'd20794, 16'd18065, 16'd62896, 16'd28985}; // indx = 4065
    #10;
    addra = 32'd130112;
    dina = {96'd0, 16'd62818, 16'd23201, 16'd8519, 16'd26769, 16'd59285, 16'd30714, 16'd35054, 16'd14161, 16'd31376, 16'd32941}; // indx = 4066
    #10;
    addra = 32'd130144;
    dina = {96'd0, 16'd50363, 16'd46315, 16'd32133, 16'd37353, 16'd34737, 16'd51386, 16'd61140, 16'd17151, 16'd44095, 16'd43098}; // indx = 4067
    #10;
    addra = 32'd130176;
    dina = {96'd0, 16'd27450, 16'd27724, 16'd25554, 16'd22833, 16'd2010, 16'd55567, 16'd43866, 16'd8486, 16'd36278, 16'd41947}; // indx = 4068
    #10;
    addra = 32'd130208;
    dina = {96'd0, 16'd13824, 16'd14300, 16'd27633, 16'd51424, 16'd3046, 16'd21086, 16'd58765, 16'd46316, 16'd23092, 16'd2044}; // indx = 4069
    #10;
    addra = 32'd130240;
    dina = {96'd0, 16'd3312, 16'd60551, 16'd16306, 16'd29289, 16'd32390, 16'd23465, 16'd36442, 16'd15193, 16'd43055, 16'd58562}; // indx = 4070
    #10;
    addra = 32'd130272;
    dina = {96'd0, 16'd64738, 16'd25052, 16'd40886, 16'd9359, 16'd34228, 16'd46704, 16'd30391, 16'd38289, 16'd51681, 16'd63070}; // indx = 4071
    #10;
    addra = 32'd130304;
    dina = {96'd0, 16'd19755, 16'd29107, 16'd49799, 16'd62302, 16'd12784, 16'd64837, 16'd11712, 16'd35031, 16'd35838, 16'd18546}; // indx = 4072
    #10;
    addra = 32'd130336;
    dina = {96'd0, 16'd22678, 16'd21920, 16'd59596, 16'd37288, 16'd970, 16'd50275, 16'd50141, 16'd32931, 16'd36377, 16'd12344}; // indx = 4073
    #10;
    addra = 32'd130368;
    dina = {96'd0, 16'd1118, 16'd43294, 16'd57357, 16'd60199, 16'd20607, 16'd22642, 16'd28062, 16'd33495, 16'd1504, 16'd30083}; // indx = 4074
    #10;
    addra = 32'd130400;
    dina = {96'd0, 16'd49571, 16'd42765, 16'd43993, 16'd54311, 16'd24015, 16'd51674, 16'd23130, 16'd24306, 16'd51295, 16'd16491}; // indx = 4075
    #10;
    addra = 32'd130432;
    dina = {96'd0, 16'd28952, 16'd3662, 16'd352, 16'd27385, 16'd1912, 16'd48323, 16'd14866, 16'd62431, 16'd43058, 16'd40929}; // indx = 4076
    #10;
    addra = 32'd130464;
    dina = {96'd0, 16'd52110, 16'd51791, 16'd14148, 16'd4058, 16'd44985, 16'd10318, 16'd38106, 16'd35324, 16'd51825, 16'd33945}; // indx = 4077
    #10;
    addra = 32'd130496;
    dina = {96'd0, 16'd16835, 16'd12471, 16'd26319, 16'd56325, 16'd30228, 16'd56316, 16'd29710, 16'd36876, 16'd19868, 16'd2935}; // indx = 4078
    #10;
    addra = 32'd130528;
    dina = {96'd0, 16'd58093, 16'd50120, 16'd53077, 16'd46040, 16'd34644, 16'd25523, 16'd20122, 16'd64393, 16'd13098, 16'd51349}; // indx = 4079
    #10;
    addra = 32'd130560;
    dina = {96'd0, 16'd54761, 16'd45880, 16'd61762, 16'd37330, 16'd31385, 16'd33246, 16'd34608, 16'd54784, 16'd47207, 16'd25226}; // indx = 4080
    #10;
    addra = 32'd130592;
    dina = {96'd0, 16'd20225, 16'd2413, 16'd31179, 16'd47105, 16'd42765, 16'd40934, 16'd36255, 16'd23425, 16'd5006, 16'd45605}; // indx = 4081
    #10;
    addra = 32'd130624;
    dina = {96'd0, 16'd20936, 16'd59750, 16'd24569, 16'd13309, 16'd54989, 16'd56718, 16'd47896, 16'd57060, 16'd1691, 16'd57258}; // indx = 4082
    #10;
    addra = 32'd130656;
    dina = {96'd0, 16'd29843, 16'd6145, 16'd46140, 16'd20531, 16'd27882, 16'd21748, 16'd23097, 16'd22625, 16'd51961, 16'd20579}; // indx = 4083
    #10;
    addra = 32'd130688;
    dina = {96'd0, 16'd53127, 16'd59713, 16'd63837, 16'd12170, 16'd32876, 16'd81, 16'd30502, 16'd7882, 16'd33899, 16'd21480}; // indx = 4084
    #10;
    addra = 32'd130720;
    dina = {96'd0, 16'd50355, 16'd14517, 16'd57957, 16'd8942, 16'd12619, 16'd63727, 16'd33470, 16'd64252, 16'd46136, 16'd36527}; // indx = 4085
    #10;
    addra = 32'd130752;
    dina = {96'd0, 16'd13939, 16'd35070, 16'd46122, 16'd18297, 16'd32848, 16'd17695, 16'd41382, 16'd20061, 16'd57928, 16'd6439}; // indx = 4086
    #10;
    addra = 32'd130784;
    dina = {96'd0, 16'd4167, 16'd16595, 16'd59703, 16'd5922, 16'd47982, 16'd47791, 16'd9620, 16'd56262, 16'd14483, 16'd51779}; // indx = 4087
    #10;
    addra = 32'd130816;
    dina = {96'd0, 16'd52995, 16'd44157, 16'd2675, 16'd12172, 16'd42650, 16'd57000, 16'd13917, 16'd51647, 16'd14645, 16'd49669}; // indx = 4088
    #10;
    addra = 32'd130848;
    dina = {96'd0, 16'd22295, 16'd23549, 16'd12471, 16'd21270, 16'd23399, 16'd48658, 16'd28946, 16'd59044, 16'd30642, 16'd64213}; // indx = 4089
    #10;
    addra = 32'd130880;
    dina = {96'd0, 16'd47515, 16'd55017, 16'd25310, 16'd2300, 16'd55637, 16'd50450, 16'd53139, 16'd12980, 16'd36208, 16'd38419}; // indx = 4090
    #10;
    addra = 32'd130912;
    dina = {96'd0, 16'd28619, 16'd21764, 16'd2327, 16'd42721, 16'd18405, 16'd64814, 16'd12319, 16'd8277, 16'd446, 16'd1920}; // indx = 4091
    #10;
    addra = 32'd130944;
    dina = {96'd0, 16'd58653, 16'd16896, 16'd42534, 16'd58965, 16'd52704, 16'd35485, 16'd13601, 16'd50697, 16'd10558, 16'd15918}; // indx = 4092
    #10;
    addra = 32'd130976;
    dina = {96'd0, 16'd50272, 16'd41367, 16'd45753, 16'd54947, 16'd55121, 16'd59017, 16'd7160, 16'd21347, 16'd4976, 16'd60494}; // indx = 4093
    #10;
    addra = 32'd131008;
    dina = {96'd0, 16'd62681, 16'd35939, 16'd12326, 16'd55033, 16'd52140, 16'd615, 16'd27593, 16'd8335, 16'd47026, 16'd2980}; // indx = 4094
    #10;
    addra = 32'd131040;
    dina = {96'd0, 16'd44860, 16'd61656, 16'd8102, 16'd63315, 16'd21897, 16'd12429, 16'd60487, 16'd38428, 16'd5728, 16'd12639}; // indx = 4095
    #10;
    addra = 32'd131072;
    dina = {96'd0, 16'd56021, 16'd40659, 16'd4397, 16'd20660, 16'd47469, 16'd25028, 16'd2761, 16'd15740, 16'd25194, 16'd9343}; // indx = 4096
    #10;
    addra = 32'd131104;
    dina = {96'd0, 16'd22915, 16'd52622, 16'd38685, 16'd55618, 16'd58308, 16'd39007, 16'd18329, 16'd55087, 16'd59809, 16'd7698}; // indx = 4097
    #10;
    addra = 32'd131136;
    dina = {96'd0, 16'd6336, 16'd54361, 16'd43752, 16'd45013, 16'd54404, 16'd39184, 16'd58403, 16'd30374, 16'd3240, 16'd23716}; // indx = 4098
    #10;
    addra = 32'd131168;
    dina = {96'd0, 16'd6015, 16'd15853, 16'd29417, 16'd15391, 16'd46227, 16'd39948, 16'd59459, 16'd26737, 16'd51723, 16'd55626}; // indx = 4099
    #10;
    addra = 32'd131200;
    dina = {96'd0, 16'd25633, 16'd7880, 16'd39184, 16'd19322, 16'd10005, 16'd1066, 16'd16763, 16'd21957, 16'd25264, 16'd16696}; // indx = 4100
    #10;
    addra = 32'd131232;
    dina = {96'd0, 16'd32177, 16'd1406, 16'd13660, 16'd48084, 16'd15001, 16'd51650, 16'd7137, 16'd14955, 16'd35160, 16'd36984}; // indx = 4101
    #10;
    addra = 32'd131264;
    dina = {96'd0, 16'd59075, 16'd42345, 16'd55913, 16'd39547, 16'd49754, 16'd30218, 16'd60200, 16'd40160, 16'd56673, 16'd717}; // indx = 4102
    #10;
    addra = 32'd131296;
    dina = {96'd0, 16'd35618, 16'd60618, 16'd18526, 16'd2462, 16'd40962, 16'd23726, 16'd4059, 16'd34210, 16'd50089, 16'd15947}; // indx = 4103
    #10;
    addra = 32'd131328;
    dina = {96'd0, 16'd23330, 16'd51496, 16'd34796, 16'd55206, 16'd48885, 16'd29429, 16'd61197, 16'd63112, 16'd13102, 16'd17474}; // indx = 4104
    #10;
    addra = 32'd131360;
    dina = {96'd0, 16'd9219, 16'd37198, 16'd20090, 16'd35102, 16'd48627, 16'd48275, 16'd31825, 16'd9187, 16'd408, 16'd54237}; // indx = 4105
    #10;
    addra = 32'd131392;
    dina = {96'd0, 16'd2315, 16'd4704, 16'd55150, 16'd43819, 16'd38143, 16'd12270, 16'd17925, 16'd46499, 16'd63471, 16'd42298}; // indx = 4106
    #10;
    addra = 32'd131424;
    dina = {96'd0, 16'd48251, 16'd2084, 16'd26029, 16'd16256, 16'd5062, 16'd49477, 16'd65023, 16'd7513, 16'd49646, 16'd47721}; // indx = 4107
    #10;
    addra = 32'd131456;
    dina = {96'd0, 16'd63639, 16'd9178, 16'd43277, 16'd34461, 16'd61676, 16'd64899, 16'd3497, 16'd45645, 16'd18442, 16'd63749}; // indx = 4108
    #10;
    addra = 32'd131488;
    dina = {96'd0, 16'd44368, 16'd7519, 16'd25638, 16'd57525, 16'd61846, 16'd9331, 16'd2502, 16'd58343, 16'd4050, 16'd25753}; // indx = 4109
    #10;
    addra = 32'd131520;
    dina = {96'd0, 16'd5301, 16'd46555, 16'd40172, 16'd11963, 16'd47522, 16'd46115, 16'd61394, 16'd40322, 16'd54142, 16'd53781}; // indx = 4110
    #10;
    addra = 32'd131552;
    dina = {96'd0, 16'd49607, 16'd26124, 16'd59336, 16'd28235, 16'd53395, 16'd44044, 16'd65036, 16'd3133, 16'd35023, 16'd16733}; // indx = 4111
    #10;
    addra = 32'd131584;
    dina = {96'd0, 16'd2065, 16'd22163, 16'd61543, 16'd16371, 16'd29412, 16'd65083, 16'd5610, 16'd342, 16'd23968, 16'd30626}; // indx = 4112
    #10;
    addra = 32'd131616;
    dina = {96'd0, 16'd15984, 16'd63837, 16'd24832, 16'd19360, 16'd30898, 16'd26275, 16'd60535, 16'd44449, 16'd18366, 16'd36894}; // indx = 4113
    #10;
    addra = 32'd131648;
    dina = {96'd0, 16'd58248, 16'd39215, 16'd46199, 16'd50376, 16'd45191, 16'd14832, 16'd14920, 16'd37500, 16'd54725, 16'd64900}; // indx = 4114
    #10;
    addra = 32'd131680;
    dina = {96'd0, 16'd7487, 16'd16531, 16'd22406, 16'd15537, 16'd24504, 16'd31365, 16'd36762, 16'd26051, 16'd49503, 16'd4822}; // indx = 4115
    #10;
    addra = 32'd131712;
    dina = {96'd0, 16'd32586, 16'd49402, 16'd20117, 16'd62238, 16'd10060, 16'd34294, 16'd4471, 16'd23307, 16'd19650, 16'd34165}; // indx = 4116
    #10;
    addra = 32'd131744;
    dina = {96'd0, 16'd16639, 16'd65278, 16'd12327, 16'd54594, 16'd22278, 16'd1985, 16'd22553, 16'd45360, 16'd62608, 16'd47007}; // indx = 4117
    #10;
    addra = 32'd131776;
    dina = {96'd0, 16'd62754, 16'd5725, 16'd28551, 16'd14302, 16'd496, 16'd35048, 16'd56223, 16'd35830, 16'd42940, 16'd49773}; // indx = 4118
    #10;
    addra = 32'd131808;
    dina = {96'd0, 16'd2937, 16'd37349, 16'd29437, 16'd51006, 16'd9574, 16'd30787, 16'd47644, 16'd56253, 16'd50552, 16'd29363}; // indx = 4119
    #10;
    addra = 32'd131840;
    dina = {96'd0, 16'd38367, 16'd57709, 16'd51168, 16'd12257, 16'd43490, 16'd54539, 16'd1456, 16'd45468, 16'd42543, 16'd2069}; // indx = 4120
    #10;
    addra = 32'd131872;
    dina = {96'd0, 16'd30235, 16'd64170, 16'd58770, 16'd29143, 16'd8263, 16'd7596, 16'd11265, 16'd21169, 16'd52618, 16'd25486}; // indx = 4121
    #10;
    addra = 32'd131904;
    dina = {96'd0, 16'd58754, 16'd54111, 16'd20096, 16'd25815, 16'd21711, 16'd53697, 16'd29310, 16'd5971, 16'd19916, 16'd45826}; // indx = 4122
    #10;
    addra = 32'd131936;
    dina = {96'd0, 16'd47131, 16'd13956, 16'd8045, 16'd30198, 16'd44883, 16'd37366, 16'd29889, 16'd57317, 16'd44454, 16'd42363}; // indx = 4123
    #10;
    addra = 32'd131968;
    dina = {96'd0, 16'd14926, 16'd22374, 16'd27743, 16'd36798, 16'd16808, 16'd56862, 16'd36851, 16'd28831, 16'd65102, 16'd9815}; // indx = 4124
    #10;
    addra = 32'd132000;
    dina = {96'd0, 16'd52887, 16'd16728, 16'd30794, 16'd6208, 16'd19588, 16'd10181, 16'd18927, 16'd40844, 16'd64947, 16'd5497}; // indx = 4125
    #10;
    addra = 32'd132032;
    dina = {96'd0, 16'd20178, 16'd10215, 16'd50195, 16'd58676, 16'd27832, 16'd46700, 16'd13533, 16'd51708, 16'd2432, 16'd23379}; // indx = 4126
    #10;
    addra = 32'd132064;
    dina = {96'd0, 16'd12640, 16'd17416, 16'd20562, 16'd30982, 16'd43569, 16'd27349, 16'd17000, 16'd15201, 16'd7874, 16'd42817}; // indx = 4127
    #10;
    addra = 32'd132096;
    dina = {96'd0, 16'd6812, 16'd22484, 16'd32608, 16'd52156, 16'd30495, 16'd26638, 16'd22946, 16'd22815, 16'd11206, 16'd36747}; // indx = 4128
    #10;
    addra = 32'd132128;
    dina = {96'd0, 16'd8712, 16'd64961, 16'd58632, 16'd14469, 16'd64921, 16'd43534, 16'd54970, 16'd45157, 16'd52245, 16'd55020}; // indx = 4129
    #10;
    addra = 32'd132160;
    dina = {96'd0, 16'd47932, 16'd52074, 16'd56014, 16'd27290, 16'd42273, 16'd30253, 16'd32435, 16'd2710, 16'd43895, 16'd25560}; // indx = 4130
    #10;
    addra = 32'd132192;
    dina = {96'd0, 16'd36380, 16'd17807, 16'd42717, 16'd6858, 16'd37871, 16'd27872, 16'd47516, 16'd28641, 16'd14435, 16'd19970}; // indx = 4131
    #10;
    addra = 32'd132224;
    dina = {96'd0, 16'd27712, 16'd23820, 16'd55369, 16'd205, 16'd23871, 16'd13011, 16'd28591, 16'd39993, 16'd36380, 16'd57436}; // indx = 4132
    #10;
    addra = 32'd132256;
    dina = {96'd0, 16'd52006, 16'd22807, 16'd33078, 16'd18697, 16'd64802, 16'd16220, 16'd1531, 16'd52802, 16'd6783, 16'd43364}; // indx = 4133
    #10;
    addra = 32'd132288;
    dina = {96'd0, 16'd50378, 16'd63841, 16'd50027, 16'd42496, 16'd58103, 16'd640, 16'd55118, 16'd29332, 16'd11926, 16'd54379}; // indx = 4134
    #10;
    addra = 32'd132320;
    dina = {96'd0, 16'd29369, 16'd40701, 16'd29137, 16'd21026, 16'd17023, 16'd37073, 16'd18940, 16'd62076, 16'd47245, 16'd15113}; // indx = 4135
    #10;
    addra = 32'd132352;
    dina = {96'd0, 16'd8056, 16'd64139, 16'd19741, 16'd57471, 16'd20511, 16'd34519, 16'd39627, 16'd33476, 16'd61074, 16'd52528}; // indx = 4136
    #10;
    addra = 32'd132384;
    dina = {96'd0, 16'd24596, 16'd39542, 16'd63963, 16'd38323, 16'd18461, 16'd12624, 16'd64132, 16'd24087, 16'd5269, 16'd38421}; // indx = 4137
    #10;
    addra = 32'd132416;
    dina = {96'd0, 16'd8720, 16'd5610, 16'd61962, 16'd22478, 16'd11170, 16'd63637, 16'd40645, 16'd11998, 16'd59058, 16'd3728}; // indx = 4138
    #10;
    addra = 32'd132448;
    dina = {96'd0, 16'd56445, 16'd39784, 16'd7069, 16'd40247, 16'd53520, 16'd37747, 16'd56118, 16'd1888, 16'd49612, 16'd65197}; // indx = 4139
    #10;
    addra = 32'd132480;
    dina = {96'd0, 16'd3593, 16'd10264, 16'd35211, 16'd26925, 16'd19808, 16'd63662, 16'd59161, 16'd14906, 16'd43103, 16'd54967}; // indx = 4140
    #10;
    addra = 32'd132512;
    dina = {96'd0, 16'd15194, 16'd20917, 16'd20530, 16'd31270, 16'd459, 16'd35149, 16'd27939, 16'd45881, 16'd20479, 16'd35516}; // indx = 4141
    #10;
    addra = 32'd132544;
    dina = {96'd0, 16'd24768, 16'd62449, 16'd4692, 16'd51077, 16'd18288, 16'd60662, 16'd35760, 16'd3424, 16'd8613, 16'd50857}; // indx = 4142
    #10;
    addra = 32'd132576;
    dina = {96'd0, 16'd42531, 16'd8659, 16'd6856, 16'd1668, 16'd33915, 16'd57114, 16'd50223, 16'd7780, 16'd24232, 16'd36645}; // indx = 4143
    #10;
    addra = 32'd132608;
    dina = {96'd0, 16'd38677, 16'd14835, 16'd33992, 16'd44665, 16'd6964, 16'd2517, 16'd32782, 16'd61009, 16'd32550, 16'd24263}; // indx = 4144
    #10;
    addra = 32'd132640;
    dina = {96'd0, 16'd18303, 16'd20174, 16'd63799, 16'd30934, 16'd64641, 16'd26712, 16'd54586, 16'd54001, 16'd9477, 16'd32657}; // indx = 4145
    #10;
    addra = 32'd132672;
    dina = {96'd0, 16'd54105, 16'd10645, 16'd32738, 16'd26249, 16'd31274, 16'd25369, 16'd43692, 16'd6350, 16'd57895, 16'd16731}; // indx = 4146
    #10;
    addra = 32'd132704;
    dina = {96'd0, 16'd31902, 16'd29105, 16'd46136, 16'd50312, 16'd35142, 16'd60214, 16'd59648, 16'd30067, 16'd20839, 16'd3762}; // indx = 4147
    #10;
    addra = 32'd132736;
    dina = {96'd0, 16'd6057, 16'd14033, 16'd116, 16'd14775, 16'd40401, 16'd20024, 16'd19257, 16'd32957, 16'd51304, 16'd45794}; // indx = 4148
    #10;
    addra = 32'd132768;
    dina = {96'd0, 16'd56619, 16'd15574, 16'd31322, 16'd6696, 16'd21011, 16'd55369, 16'd8105, 16'd36268, 16'd18923, 16'd19070}; // indx = 4149
    #10;
    addra = 32'd132800;
    dina = {96'd0, 16'd47801, 16'd31852, 16'd13604, 16'd22203, 16'd39368, 16'd45947, 16'd12541, 16'd58715, 16'd53996, 16'd1245}; // indx = 4150
    #10;
    addra = 32'd132832;
    dina = {96'd0, 16'd8730, 16'd33594, 16'd16886, 16'd24628, 16'd7121, 16'd10293, 16'd46742, 16'd32945, 16'd59335, 16'd38735}; // indx = 4151
    #10;
    addra = 32'd132864;
    dina = {96'd0, 16'd2289, 16'd22390, 16'd12650, 16'd20880, 16'd11550, 16'd9241, 16'd60050, 16'd18684, 16'd47170, 16'd23493}; // indx = 4152
    #10;
    addra = 32'd132896;
    dina = {96'd0, 16'd65187, 16'd8829, 16'd59881, 16'd1054, 16'd27831, 16'd12236, 16'd20618, 16'd2530, 16'd42875, 16'd40017}; // indx = 4153
    #10;
    addra = 32'd132928;
    dina = {96'd0, 16'd29971, 16'd42606, 16'd14412, 16'd39774, 16'd33766, 16'd1378, 16'd37485, 16'd41514, 16'd38448, 16'd11670}; // indx = 4154
    #10;
    addra = 32'd132960;
    dina = {96'd0, 16'd38556, 16'd44308, 16'd23902, 16'd13917, 16'd17537, 16'd6384, 16'd24985, 16'd20876, 16'd7792, 16'd21507}; // indx = 4155
    #10;
    addra = 32'd132992;
    dina = {96'd0, 16'd40286, 16'd61268, 16'd18076, 16'd7103, 16'd47318, 16'd16559, 16'd38053, 16'd3418, 16'd44440, 16'd17190}; // indx = 4156
    #10;
    addra = 32'd133024;
    dina = {96'd0, 16'd36442, 16'd40641, 16'd30771, 16'd33555, 16'd34572, 16'd39350, 16'd51160, 16'd219, 16'd61147, 16'd43357}; // indx = 4157
    #10;
    addra = 32'd133056;
    dina = {96'd0, 16'd38925, 16'd31888, 16'd25974, 16'd1260, 16'd29657, 16'd42613, 16'd57750, 16'd4876, 16'd13855, 16'd6784}; // indx = 4158
    #10;
    addra = 32'd133088;
    dina = {96'd0, 16'd52811, 16'd32691, 16'd40427, 16'd14212, 16'd2362, 16'd15314, 16'd28427, 16'd53664, 16'd9376, 16'd42148}; // indx = 4159
    #10;
    addra = 32'd133120;
    dina = {96'd0, 16'd47958, 16'd45548, 16'd58887, 16'd64677, 16'd14261, 16'd29534, 16'd57604, 16'd55036, 16'd36664, 16'd14257}; // indx = 4160
    #10;
    addra = 32'd133152;
    dina = {96'd0, 16'd6102, 16'd32681, 16'd13145, 16'd25989, 16'd55605, 16'd54736, 16'd6147, 16'd33215, 16'd50449, 16'd63882}; // indx = 4161
    #10;
    addra = 32'd133184;
    dina = {96'd0, 16'd62649, 16'd11563, 16'd25446, 16'd33226, 16'd37999, 16'd38600, 16'd6587, 16'd40615, 16'd20082, 16'd33153}; // indx = 4162
    #10;
    addra = 32'd133216;
    dina = {96'd0, 16'd4074, 16'd16463, 16'd10046, 16'd55155, 16'd25841, 16'd38728, 16'd46206, 16'd3105, 16'd5957, 16'd46575}; // indx = 4163
    #10;
    addra = 32'd133248;
    dina = {96'd0, 16'd4776, 16'd8889, 16'd36961, 16'd1342, 16'd38987, 16'd41968, 16'd29664, 16'd33408, 16'd62917, 16'd19274}; // indx = 4164
    #10;
    addra = 32'd133280;
    dina = {96'd0, 16'd692, 16'd11306, 16'd7031, 16'd53148, 16'd41010, 16'd26798, 16'd38739, 16'd1201, 16'd27824, 16'd13554}; // indx = 4165
    #10;
    addra = 32'd133312;
    dina = {96'd0, 16'd47343, 16'd14419, 16'd19634, 16'd10445, 16'd6267, 16'd2483, 16'd47176, 16'd866, 16'd17962, 16'd10148}; // indx = 4166
    #10;
    addra = 32'd133344;
    dina = {96'd0, 16'd43829, 16'd12069, 16'd24825, 16'd34610, 16'd38503, 16'd16520, 16'd46398, 16'd62008, 16'd6530, 16'd40482}; // indx = 4167
    #10;
    addra = 32'd133376;
    dina = {96'd0, 16'd9973, 16'd40325, 16'd62860, 16'd64081, 16'd51453, 16'd44147, 16'd49618, 16'd43390, 16'd31861, 16'd7993}; // indx = 4168
    #10;
    addra = 32'd133408;
    dina = {96'd0, 16'd52108, 16'd12182, 16'd56136, 16'd48579, 16'd59094, 16'd35139, 16'd55158, 16'd23433, 16'd16515, 16'd30464}; // indx = 4169
    #10;
    addra = 32'd133440;
    dina = {96'd0, 16'd1534, 16'd46736, 16'd33011, 16'd36114, 16'd473, 16'd63095, 16'd57148, 16'd26792, 16'd45046, 16'd13398}; // indx = 4170
    #10;
    addra = 32'd133472;
    dina = {96'd0, 16'd42084, 16'd17429, 16'd41141, 16'd17498, 16'd63948, 16'd45948, 16'd15980, 16'd21295, 16'd64274, 16'd33899}; // indx = 4171
    #10;
    addra = 32'd133504;
    dina = {96'd0, 16'd55344, 16'd17253, 16'd22565, 16'd28011, 16'd54078, 16'd38286, 16'd6658, 16'd42153, 16'd18166, 16'd24900}; // indx = 4172
    #10;
    addra = 32'd133536;
    dina = {96'd0, 16'd42180, 16'd55705, 16'd39307, 16'd11118, 16'd64377, 16'd47557, 16'd59947, 16'd1896, 16'd18933, 16'd26075}; // indx = 4173
    #10;
    addra = 32'd133568;
    dina = {96'd0, 16'd29871, 16'd17325, 16'd62280, 16'd32333, 16'd2540, 16'd53460, 16'd59021, 16'd37962, 16'd33008, 16'd50263}; // indx = 4174
    #10;
    addra = 32'd133600;
    dina = {96'd0, 16'd8745, 16'd27639, 16'd41085, 16'd29374, 16'd17341, 16'd42852, 16'd14043, 16'd52453, 16'd44986, 16'd10516}; // indx = 4175
    #10;
    addra = 32'd133632;
    dina = {96'd0, 16'd13555, 16'd42299, 16'd30965, 16'd23314, 16'd30564, 16'd43784, 16'd47051, 16'd29082, 16'd14018, 16'd8632}; // indx = 4176
    #10;
    addra = 32'd133664;
    dina = {96'd0, 16'd51276, 16'd39868, 16'd11164, 16'd51918, 16'd40278, 16'd37557, 16'd41232, 16'd26750, 16'd29751, 16'd15215}; // indx = 4177
    #10;
    addra = 32'd133696;
    dina = {96'd0, 16'd27073, 16'd63632, 16'd35870, 16'd57219, 16'd58695, 16'd27669, 16'd4744, 16'd34886, 16'd50458, 16'd58675}; // indx = 4178
    #10;
    addra = 32'd133728;
    dina = {96'd0, 16'd4984, 16'd54881, 16'd64929, 16'd37337, 16'd65156, 16'd57511, 16'd33296, 16'd62961, 16'd30539, 16'd33470}; // indx = 4179
    #10;
    addra = 32'd133760;
    dina = {96'd0, 16'd55541, 16'd46872, 16'd59809, 16'd59035, 16'd58201, 16'd23668, 16'd27351, 16'd32531, 16'd45947, 16'd744}; // indx = 4180
    #10;
    addra = 32'd133792;
    dina = {96'd0, 16'd48445, 16'd32416, 16'd32894, 16'd21996, 16'd27196, 16'd9222, 16'd52546, 16'd11202, 16'd36048, 16'd48078}; // indx = 4181
    #10;
    addra = 32'd133824;
    dina = {96'd0, 16'd39641, 16'd33773, 16'd18239, 16'd60581, 16'd54955, 16'd46380, 16'd37834, 16'd35874, 16'd2458, 16'd12898}; // indx = 4182
    #10;
    addra = 32'd133856;
    dina = {96'd0, 16'd50571, 16'd48516, 16'd12707, 16'd2081, 16'd17841, 16'd5391, 16'd36639, 16'd64987, 16'd36092, 16'd56207}; // indx = 4183
    #10;
    addra = 32'd133888;
    dina = {96'd0, 16'd1723, 16'd25197, 16'd54115, 16'd46726, 16'd26586, 16'd6599, 16'd45039, 16'd56118, 16'd14697, 16'd55627}; // indx = 4184
    #10;
    addra = 32'd133920;
    dina = {96'd0, 16'd14579, 16'd8702, 16'd37860, 16'd22125, 16'd58688, 16'd56031, 16'd63169, 16'd5919, 16'd45857, 16'd13336}; // indx = 4185
    #10;
    addra = 32'd133952;
    dina = {96'd0, 16'd19820, 16'd46628, 16'd42523, 16'd50520, 16'd30581, 16'd24773, 16'd18504, 16'd47269, 16'd60319, 16'd64580}; // indx = 4186
    #10;
    addra = 32'd133984;
    dina = {96'd0, 16'd53353, 16'd56612, 16'd57860, 16'd36301, 16'd14442, 16'd28789, 16'd10708, 16'd47781, 16'd26014, 16'd31681}; // indx = 4187
    #10;
    addra = 32'd134016;
    dina = {96'd0, 16'd14237, 16'd21252, 16'd25875, 16'd45152, 16'd10295, 16'd36564, 16'd15509, 16'd36290, 16'd26134, 16'd10642}; // indx = 4188
    #10;
    addra = 32'd134048;
    dina = {96'd0, 16'd20327, 16'd16439, 16'd27283, 16'd29308, 16'd36084, 16'd64238, 16'd41024, 16'd3655, 16'd1227, 16'd54639}; // indx = 4189
    #10;
    addra = 32'd134080;
    dina = {96'd0, 16'd33882, 16'd13631, 16'd50724, 16'd35414, 16'd18680, 16'd9933, 16'd39245, 16'd32398, 16'd37272, 16'd8508}; // indx = 4190
    #10;
    addra = 32'd134112;
    dina = {96'd0, 16'd19436, 16'd33950, 16'd39540, 16'd14856, 16'd54237, 16'd6501, 16'd32347, 16'd18604, 16'd41019, 16'd17772}; // indx = 4191
    #10;
    addra = 32'd134144;
    dina = {96'd0, 16'd4727, 16'd28778, 16'd23530, 16'd507, 16'd27659, 16'd34576, 16'd56716, 16'd34753, 16'd39745, 16'd26571}; // indx = 4192
    #10;
    addra = 32'd134176;
    dina = {96'd0, 16'd43091, 16'd32108, 16'd2884, 16'd3707, 16'd57761, 16'd5277, 16'd40816, 16'd35595, 16'd12732, 16'd1980}; // indx = 4193
    #10;
    addra = 32'd134208;
    dina = {96'd0, 16'd37412, 16'd42044, 16'd21172, 16'd24305, 16'd7582, 16'd9429, 16'd6790, 16'd21600, 16'd37193, 16'd1482}; // indx = 4194
    #10;
    addra = 32'd134240;
    dina = {96'd0, 16'd49119, 16'd9449, 16'd34052, 16'd57202, 16'd26705, 16'd64661, 16'd41435, 16'd6582, 16'd37351, 16'd64323}; // indx = 4195
    #10;
    addra = 32'd134272;
    dina = {96'd0, 16'd44777, 16'd4662, 16'd46241, 16'd10834, 16'd441, 16'd48519, 16'd57238, 16'd3566, 16'd58774, 16'd18452}; // indx = 4196
    #10;
    addra = 32'd134304;
    dina = {96'd0, 16'd19913, 16'd11969, 16'd60313, 16'd3793, 16'd1826, 16'd40850, 16'd16518, 16'd13416, 16'd28317, 16'd55103}; // indx = 4197
    #10;
    addra = 32'd134336;
    dina = {96'd0, 16'd40326, 16'd33456, 16'd46457, 16'd65003, 16'd42806, 16'd50836, 16'd58560, 16'd26420, 16'd11637, 16'd7938}; // indx = 4198
    #10;
    addra = 32'd134368;
    dina = {96'd0, 16'd46386, 16'd44102, 16'd15228, 16'd26596, 16'd30324, 16'd45015, 16'd61289, 16'd60793, 16'd38926, 16'd33468}; // indx = 4199
    #10;
    addra = 32'd134400;
    dina = {96'd0, 16'd17557, 16'd46275, 16'd31923, 16'd28890, 16'd26764, 16'd64764, 16'd18409, 16'd8293, 16'd33637, 16'd26120}; // indx = 4200
    #10;
    addra = 32'd134432;
    dina = {96'd0, 16'd54820, 16'd25608, 16'd49852, 16'd51515, 16'd1192, 16'd18814, 16'd32698, 16'd35552, 16'd9123, 16'd1194}; // indx = 4201
    #10;
    addra = 32'd134464;
    dina = {96'd0, 16'd63022, 16'd45624, 16'd18523, 16'd414, 16'd52916, 16'd56168, 16'd50789, 16'd44624, 16'd36780, 16'd17012}; // indx = 4202
    #10;
    addra = 32'd134496;
    dina = {96'd0, 16'd28103, 16'd22363, 16'd6025, 16'd51596, 16'd31510, 16'd44445, 16'd24965, 16'd25480, 16'd18875, 16'd25151}; // indx = 4203
    #10;
    addra = 32'd134528;
    dina = {96'd0, 16'd1284, 16'd62875, 16'd22719, 16'd64391, 16'd8122, 16'd11005, 16'd61555, 16'd18343, 16'd3924, 16'd63081}; // indx = 4204
    #10;
    addra = 32'd134560;
    dina = {96'd0, 16'd44638, 16'd7208, 16'd27937, 16'd32204, 16'd38603, 16'd18083, 16'd56679, 16'd43362, 16'd43554, 16'd17291}; // indx = 4205
    #10;
    addra = 32'd134592;
    dina = {96'd0, 16'd34982, 16'd18469, 16'd7312, 16'd14552, 16'd34970, 16'd42560, 16'd19064, 16'd22316, 16'd39976, 16'd41558}; // indx = 4206
    #10;
    addra = 32'd134624;
    dina = {96'd0, 16'd49457, 16'd30692, 16'd31568, 16'd23050, 16'd37146, 16'd11685, 16'd16124, 16'd57374, 16'd46263, 16'd30312}; // indx = 4207
    #10;
    addra = 32'd134656;
    dina = {96'd0, 16'd14106, 16'd44916, 16'd7934, 16'd55179, 16'd1448, 16'd1002, 16'd37627, 16'd40299, 16'd63532, 16'd27460}; // indx = 4208
    #10;
    addra = 32'd134688;
    dina = {96'd0, 16'd23153, 16'd61923, 16'd17427, 16'd58037, 16'd39817, 16'd38739, 16'd31187, 16'd20365, 16'd19382, 16'd57315}; // indx = 4209
    #10;
    addra = 32'd134720;
    dina = {96'd0, 16'd65352, 16'd51791, 16'd56283, 16'd10959, 16'd6924, 16'd16647, 16'd3061, 16'd64121, 16'd23511, 16'd51564}; // indx = 4210
    #10;
    addra = 32'd134752;
    dina = {96'd0, 16'd10319, 16'd54576, 16'd36462, 16'd13740, 16'd37770, 16'd601, 16'd15754, 16'd23951, 16'd57431, 16'd38406}; // indx = 4211
    #10;
    addra = 32'd134784;
    dina = {96'd0, 16'd20291, 16'd272, 16'd16025, 16'd35346, 16'd1577, 16'd40706, 16'd58501, 16'd43581, 16'd14772, 16'd54620}; // indx = 4212
    #10;
    addra = 32'd134816;
    dina = {96'd0, 16'd48590, 16'd30326, 16'd51911, 16'd61102, 16'd17027, 16'd24629, 16'd29879, 16'd60172, 16'd25959, 16'd51563}; // indx = 4213
    #10;
    addra = 32'd134848;
    dina = {96'd0, 16'd4287, 16'd18464, 16'd30900, 16'd55122, 16'd23077, 16'd43239, 16'd32089, 16'd29097, 16'd15340, 16'd50953}; // indx = 4214
    #10;
    addra = 32'd134880;
    dina = {96'd0, 16'd24113, 16'd47635, 16'd47089, 16'd53801, 16'd9735, 16'd16313, 16'd25193, 16'd18388, 16'd20032, 16'd55785}; // indx = 4215
    #10;
    addra = 32'd134912;
    dina = {96'd0, 16'd52707, 16'd1625, 16'd31786, 16'd18952, 16'd37894, 16'd50922, 16'd40795, 16'd31163, 16'd9848, 16'd43524}; // indx = 4216
    #10;
    addra = 32'd134944;
    dina = {96'd0, 16'd40792, 16'd20050, 16'd4081, 16'd17896, 16'd60764, 16'd25750, 16'd48599, 16'd46578, 16'd64992, 16'd5324}; // indx = 4217
    #10;
    addra = 32'd134976;
    dina = {96'd0, 16'd40118, 16'd10196, 16'd6222, 16'd31773, 16'd25296, 16'd30634, 16'd17778, 16'd60628, 16'd21290, 16'd57670}; // indx = 4218
    #10;
    addra = 32'd135008;
    dina = {96'd0, 16'd49306, 16'd64435, 16'd22079, 16'd23755, 16'd928, 16'd31908, 16'd37692, 16'd22698, 16'd40669, 16'd17893}; // indx = 4219
    #10;
    addra = 32'd135040;
    dina = {96'd0, 16'd45202, 16'd48927, 16'd55977, 16'd1872, 16'd24788, 16'd3280, 16'd53911, 16'd48582, 16'd49727, 16'd5956}; // indx = 4220
    #10;
    addra = 32'd135072;
    dina = {96'd0, 16'd36200, 16'd34999, 16'd56173, 16'd57948, 16'd27128, 16'd10370, 16'd34058, 16'd16401, 16'd4107, 16'd38233}; // indx = 4221
    #10;
    addra = 32'd135104;
    dina = {96'd0, 16'd594, 16'd24344, 16'd32283, 16'd60005, 16'd25075, 16'd39523, 16'd55677, 16'd51877, 16'd26269, 16'd6969}; // indx = 4222
    #10;
    addra = 32'd135136;
    dina = {96'd0, 16'd60475, 16'd49878, 16'd8170, 16'd1323, 16'd28719, 16'd32039, 16'd24139, 16'd48328, 16'd56439, 16'd14005}; // indx = 4223
    #10;
    addra = 32'd135168;
    dina = {96'd0, 16'd37409, 16'd59908, 16'd40531, 16'd21216, 16'd56680, 16'd54344, 16'd5355, 16'd39303, 16'd17829, 16'd41291}; // indx = 4224
    #10;
    addra = 32'd135200;
    dina = {96'd0, 16'd48907, 16'd41749, 16'd28149, 16'd791, 16'd50285, 16'd65104, 16'd39577, 16'd1374, 16'd54210, 16'd46243}; // indx = 4225
    #10;
    addra = 32'd135232;
    dina = {96'd0, 16'd63147, 16'd53449, 16'd35535, 16'd63856, 16'd53603, 16'd21427, 16'd44519, 16'd5937, 16'd59733, 16'd48718}; // indx = 4226
    #10;
    addra = 32'd135264;
    dina = {96'd0, 16'd41790, 16'd23457, 16'd4598, 16'd34611, 16'd17810, 16'd34026, 16'd63225, 16'd62802, 16'd58688, 16'd1772}; // indx = 4227
    #10;
    addra = 32'd135296;
    dina = {96'd0, 16'd3018, 16'd37546, 16'd24710, 16'd51889, 16'd35043, 16'd64635, 16'd17535, 16'd34617, 16'd39216, 16'd20113}; // indx = 4228
    #10;
    addra = 32'd135328;
    dina = {96'd0, 16'd64234, 16'd6964, 16'd2257, 16'd26057, 16'd62900, 16'd36575, 16'd60155, 16'd27221, 16'd1542, 16'd20228}; // indx = 4229
    #10;
    addra = 32'd135360;
    dina = {96'd0, 16'd60088, 16'd56873, 16'd32281, 16'd9344, 16'd50006, 16'd55089, 16'd37544, 16'd64279, 16'd41852, 16'd15112}; // indx = 4230
    #10;
    addra = 32'd135392;
    dina = {96'd0, 16'd9572, 16'd8462, 16'd45841, 16'd4693, 16'd31863, 16'd1838, 16'd27802, 16'd57888, 16'd35185, 16'd11618}; // indx = 4231
    #10;
    addra = 32'd135424;
    dina = {96'd0, 16'd42718, 16'd46971, 16'd35440, 16'd23087, 16'd47496, 16'd59512, 16'd65248, 16'd6083, 16'd4985, 16'd30240}; // indx = 4232
    #10;
    addra = 32'd135456;
    dina = {96'd0, 16'd64178, 16'd3367, 16'd267, 16'd56315, 16'd36943, 16'd21796, 16'd61460, 16'd17281, 16'd28417, 16'd29679}; // indx = 4233
    #10;
    addra = 32'd135488;
    dina = {96'd0, 16'd31416, 16'd7425, 16'd51284, 16'd51014, 16'd33456, 16'd27291, 16'd3858, 16'd11191, 16'd11578, 16'd56791}; // indx = 4234
    #10;
    addra = 32'd135520;
    dina = {96'd0, 16'd4609, 16'd31237, 16'd8707, 16'd26051, 16'd61319, 16'd12178, 16'd42501, 16'd29752, 16'd1507, 16'd13716}; // indx = 4235
    #10;
    addra = 32'd135552;
    dina = {96'd0, 16'd63830, 16'd51582, 16'd45220, 16'd45545, 16'd16073, 16'd23450, 16'd9889, 16'd26020, 16'd64608, 16'd43630}; // indx = 4236
    #10;
    addra = 32'd135584;
    dina = {96'd0, 16'd53556, 16'd18504, 16'd34629, 16'd47317, 16'd52801, 16'd19819, 16'd49870, 16'd61088, 16'd47193, 16'd21785}; // indx = 4237
    #10;
    addra = 32'd135616;
    dina = {96'd0, 16'd39096, 16'd58429, 16'd573, 16'd12482, 16'd8627, 16'd11463, 16'd19800, 16'd29954, 16'd48919, 16'd12462}; // indx = 4238
    #10;
    addra = 32'd135648;
    dina = {96'd0, 16'd54898, 16'd13456, 16'd28890, 16'd43844, 16'd3386, 16'd48126, 16'd31868, 16'd61042, 16'd52301, 16'd58392}; // indx = 4239
    #10;
    addra = 32'd135680;
    dina = {96'd0, 16'd3640, 16'd47438, 16'd4375, 16'd3232, 16'd53855, 16'd32407, 16'd53275, 16'd5720, 16'd8644, 16'd30791}; // indx = 4240
    #10;
    addra = 32'd135712;
    dina = {96'd0, 16'd15037, 16'd44343, 16'd16759, 16'd36606, 16'd57124, 16'd2457, 16'd24389, 16'd35694, 16'd37677, 16'd47591}; // indx = 4241
    #10;
    addra = 32'd135744;
    dina = {96'd0, 16'd55814, 16'd5907, 16'd32439, 16'd51359, 16'd27623, 16'd3667, 16'd64162, 16'd3938, 16'd64215, 16'd55727}; // indx = 4242
    #10;
    addra = 32'd135776;
    dina = {96'd0, 16'd42984, 16'd8262, 16'd51163, 16'd24845, 16'd65488, 16'd140, 16'd18122, 16'd32113, 16'd54199, 16'd1015}; // indx = 4243
    #10;
    addra = 32'd135808;
    dina = {96'd0, 16'd20563, 16'd58805, 16'd65535, 16'd56339, 16'd41203, 16'd39351, 16'd23953, 16'd34662, 16'd47465, 16'd15888}; // indx = 4244
    #10;
    addra = 32'd135840;
    dina = {96'd0, 16'd45194, 16'd34557, 16'd11203, 16'd35208, 16'd14259, 16'd63216, 16'd52392, 16'd50146, 16'd49913, 16'd51777}; // indx = 4245
    #10;
    addra = 32'd135872;
    dina = {96'd0, 16'd12073, 16'd31033, 16'd20830, 16'd18447, 16'd20426, 16'd24011, 16'd56844, 16'd11134, 16'd44595, 16'd35593}; // indx = 4246
    #10;
    addra = 32'd135904;
    dina = {96'd0, 16'd28537, 16'd33739, 16'd23531, 16'd24286, 16'd62402, 16'd4438, 16'd22474, 16'd21844, 16'd21959, 16'd3818}; // indx = 4247
    #10;
    addra = 32'd135936;
    dina = {96'd0, 16'd9333, 16'd61376, 16'd15268, 16'd8082, 16'd3075, 16'd261, 16'd30808, 16'd30555, 16'd62583, 16'd65453}; // indx = 4248
    #10;
    addra = 32'd135968;
    dina = {96'd0, 16'd29180, 16'd50435, 16'd53596, 16'd33106, 16'd32226, 16'd42208, 16'd48466, 16'd61351, 16'd20841, 16'd16702}; // indx = 4249
    #10;
    addra = 32'd136000;
    dina = {96'd0, 16'd40422, 16'd37711, 16'd55850, 16'd38503, 16'd51794, 16'd3604, 16'd6244, 16'd32878, 16'd10389, 16'd54122}; // indx = 4250
    #10;
    addra = 32'd136032;
    dina = {96'd0, 16'd39893, 16'd17776, 16'd10144, 16'd26502, 16'd56552, 16'd60205, 16'd13513, 16'd24238, 16'd59198, 16'd43489}; // indx = 4251
    #10;
    addra = 32'd136064;
    dina = {96'd0, 16'd3838, 16'd60510, 16'd61497, 16'd7739, 16'd33100, 16'd13505, 16'd8192, 16'd20772, 16'd8373, 16'd30963}; // indx = 4252
    #10;
    addra = 32'd136096;
    dina = {96'd0, 16'd2924, 16'd52933, 16'd44235, 16'd39453, 16'd43917, 16'd5374, 16'd32211, 16'd33556, 16'd54664, 16'd64985}; // indx = 4253
    #10;
    addra = 32'd136128;
    dina = {96'd0, 16'd61931, 16'd38295, 16'd57527, 16'd15835, 16'd64276, 16'd31914, 16'd61346, 16'd37539, 16'd58935, 16'd34120}; // indx = 4254
    #10;
    addra = 32'd136160;
    dina = {96'd0, 16'd52149, 16'd64523, 16'd32474, 16'd61119, 16'd24365, 16'd13934, 16'd52424, 16'd38636, 16'd6783, 16'd18472}; // indx = 4255
    #10;
    addra = 32'd136192;
    dina = {96'd0, 16'd51681, 16'd38702, 16'd3593, 16'd1280, 16'd39598, 16'd53629, 16'd905, 16'd30033, 16'd37719, 16'd58986}; // indx = 4256
    #10;
    addra = 32'd136224;
    dina = {96'd0, 16'd27132, 16'd15313, 16'd14370, 16'd5485, 16'd42772, 16'd12448, 16'd36783, 16'd21755, 16'd60764, 16'd45554}; // indx = 4257
    #10;
    addra = 32'd136256;
    dina = {96'd0, 16'd28859, 16'd30451, 16'd51559, 16'd16890, 16'd50956, 16'd15478, 16'd59435, 16'd9428, 16'd22464, 16'd22775}; // indx = 4258
    #10;
    addra = 32'd136288;
    dina = {96'd0, 16'd37786, 16'd49217, 16'd35760, 16'd42684, 16'd21681, 16'd32905, 16'd18789, 16'd43488, 16'd46234, 16'd11734}; // indx = 4259
    #10;
    addra = 32'd136320;
    dina = {96'd0, 16'd49967, 16'd47496, 16'd63652, 16'd39269, 16'd32302, 16'd31270, 16'd64510, 16'd34340, 16'd37902, 16'd25668}; // indx = 4260
    #10;
    addra = 32'd136352;
    dina = {96'd0, 16'd34520, 16'd9307, 16'd46258, 16'd2106, 16'd14743, 16'd24642, 16'd17424, 16'd63945, 16'd45177, 16'd24860}; // indx = 4261
    #10;
    addra = 32'd136384;
    dina = {96'd0, 16'd51917, 16'd26857, 16'd34969, 16'd24251, 16'd49380, 16'd19807, 16'd4317, 16'd43104, 16'd56106, 16'd39358}; // indx = 4262
    #10;
    addra = 32'd136416;
    dina = {96'd0, 16'd13263, 16'd14476, 16'd18067, 16'd18294, 16'd59572, 16'd17971, 16'd10515, 16'd19429, 16'd24166, 16'd62587}; // indx = 4263
    #10;
    addra = 32'd136448;
    dina = {96'd0, 16'd22937, 16'd15406, 16'd17771, 16'd58114, 16'd4315, 16'd52280, 16'd9420, 16'd23900, 16'd20173, 16'd28960}; // indx = 4264
    #10;
    addra = 32'd136480;
    dina = {96'd0, 16'd8245, 16'd49835, 16'd44581, 16'd44783, 16'd11168, 16'd30637, 16'd58357, 16'd24741, 16'd62449, 16'd32640}; // indx = 4265
    #10;
    addra = 32'd136512;
    dina = {96'd0, 16'd19423, 16'd26674, 16'd27878, 16'd64739, 16'd16478, 16'd65374, 16'd43965, 16'd6240, 16'd17317, 16'd46395}; // indx = 4266
    #10;
    addra = 32'd136544;
    dina = {96'd0, 16'd8941, 16'd61903, 16'd47189, 16'd16893, 16'd53835, 16'd38303, 16'd29569, 16'd4692, 16'd21242, 16'd12613}; // indx = 4267
    #10;
    addra = 32'd136576;
    dina = {96'd0, 16'd92, 16'd46292, 16'd49299, 16'd6499, 16'd4599, 16'd12781, 16'd63869, 16'd12423, 16'd9033, 16'd10117}; // indx = 4268
    #10;
    addra = 32'd136608;
    dina = {96'd0, 16'd1218, 16'd61574, 16'd3093, 16'd16702, 16'd25493, 16'd14639, 16'd27108, 16'd31510, 16'd13298, 16'd10655}; // indx = 4269
    #10;
    addra = 32'd136640;
    dina = {96'd0, 16'd24321, 16'd10901, 16'd55146, 16'd35307, 16'd51487, 16'd58557, 16'd10104, 16'd53072, 16'd53231, 16'd18089}; // indx = 4270
    #10;
    addra = 32'd136672;
    dina = {96'd0, 16'd36114, 16'd13380, 16'd38910, 16'd42421, 16'd641, 16'd21140, 16'd31737, 16'd38591, 16'd51681, 16'd55759}; // indx = 4271
    #10;
    addra = 32'd136704;
    dina = {96'd0, 16'd22889, 16'd48595, 16'd37112, 16'd58474, 16'd62316, 16'd39799, 16'd30860, 16'd28916, 16'd61472, 16'd38466}; // indx = 4272
    #10;
    addra = 32'd136736;
    dina = {96'd0, 16'd29123, 16'd63386, 16'd46150, 16'd55863, 16'd42636, 16'd12471, 16'd19481, 16'd22657, 16'd14446, 16'd48896}; // indx = 4273
    #10;
    addra = 32'd136768;
    dina = {96'd0, 16'd10040, 16'd34471, 16'd29481, 16'd47138, 16'd64625, 16'd57928, 16'd40857, 16'd31362, 16'd11050, 16'd28931}; // indx = 4274
    #10;
    addra = 32'd136800;
    dina = {96'd0, 16'd13441, 16'd45597, 16'd22383, 16'd59761, 16'd60502, 16'd52034, 16'd14567, 16'd3304, 16'd40661, 16'd16305}; // indx = 4275
    #10;
    addra = 32'd136832;
    dina = {96'd0, 16'd46299, 16'd56612, 16'd62720, 16'd58281, 16'd57614, 16'd2643, 16'd21110, 16'd11688, 16'd19041, 16'd22308}; // indx = 4276
    #10;
    addra = 32'd136864;
    dina = {96'd0, 16'd65498, 16'd13979, 16'd31384, 16'd42469, 16'd57639, 16'd21722, 16'd20197, 16'd3520, 16'd18411, 16'd33969}; // indx = 4277
    #10;
    addra = 32'd136896;
    dina = {96'd0, 16'd30835, 16'd42331, 16'd59955, 16'd37201, 16'd34728, 16'd48828, 16'd1575, 16'd35263, 16'd13294, 16'd55198}; // indx = 4278
    #10;
    addra = 32'd136928;
    dina = {96'd0, 16'd42936, 16'd44285, 16'd48723, 16'd37759, 16'd31505, 16'd34148, 16'd38433, 16'd59820, 16'd16649, 16'd945}; // indx = 4279
    #10;
    addra = 32'd136960;
    dina = {96'd0, 16'd16629, 16'd20502, 16'd13908, 16'd37269, 16'd8562, 16'd12276, 16'd52346, 16'd25153, 16'd47178, 16'd49054}; // indx = 4280
    #10;
    addra = 32'd136992;
    dina = {96'd0, 16'd56380, 16'd45105, 16'd44099, 16'd56270, 16'd56776, 16'd41712, 16'd53571, 16'd14947, 16'd7796, 16'd60163}; // indx = 4281
    #10;
    addra = 32'd137024;
    dina = {96'd0, 16'd8207, 16'd33332, 16'd44780, 16'd22960, 16'd28776, 16'd58679, 16'd26587, 16'd43527, 16'd18820, 16'd43065}; // indx = 4282
    #10;
    addra = 32'd137056;
    dina = {96'd0, 16'd11481, 16'd20459, 16'd8480, 16'd17712, 16'd56142, 16'd34035, 16'd25264, 16'd6220, 16'd13420, 16'd63377}; // indx = 4283
    #10;
    addra = 32'd137088;
    dina = {96'd0, 16'd35584, 16'd16266, 16'd42454, 16'd50436, 16'd16581, 16'd59358, 16'd30562, 16'd41418, 16'd31769, 16'd55524}; // indx = 4284
    #10;
    addra = 32'd137120;
    dina = {96'd0, 16'd62426, 16'd18219, 16'd2332, 16'd27939, 16'd65001, 16'd38873, 16'd64098, 16'd34563, 16'd53927, 16'd10141}; // indx = 4285
    #10;
    addra = 32'd137152;
    dina = {96'd0, 16'd4033, 16'd13024, 16'd50822, 16'd8115, 16'd51640, 16'd16068, 16'd59035, 16'd30109, 16'd32066, 16'd22928}; // indx = 4286
    #10;
    addra = 32'd137184;
    dina = {96'd0, 16'd19753, 16'd47555, 16'd59376, 16'd18896, 16'd42300, 16'd40020, 16'd47, 16'd35965, 16'd57464, 16'd50873}; // indx = 4287
    #10;
    addra = 32'd137216;
    dina = {96'd0, 16'd63572, 16'd36456, 16'd61778, 16'd27383, 16'd22065, 16'd45503, 16'd38373, 16'd24734, 16'd21235, 16'd2850}; // indx = 4288
    #10;
    addra = 32'd137248;
    dina = {96'd0, 16'd30888, 16'd46136, 16'd13761, 16'd39686, 16'd62675, 16'd36203, 16'd52488, 16'd44367, 16'd35512, 16'd16864}; // indx = 4289
    #10;
    addra = 32'd137280;
    dina = {96'd0, 16'd41750, 16'd41632, 16'd8919, 16'd13796, 16'd50152, 16'd62514, 16'd10046, 16'd44691, 16'd58148, 16'd25842}; // indx = 4290
    #10;
    addra = 32'd137312;
    dina = {96'd0, 16'd271, 16'd51489, 16'd55084, 16'd59129, 16'd62082, 16'd25776, 16'd51648, 16'd63397, 16'd63113, 16'd47376}; // indx = 4291
    #10;
    addra = 32'd137344;
    dina = {96'd0, 16'd40837, 16'd30590, 16'd24187, 16'd43610, 16'd31693, 16'd38154, 16'd1792, 16'd10176, 16'd34394, 16'd40443}; // indx = 4292
    #10;
    addra = 32'd137376;
    dina = {96'd0, 16'd57053, 16'd35178, 16'd61123, 16'd2227, 16'd19739, 16'd59832, 16'd25702, 16'd22167, 16'd46736, 16'd38700}; // indx = 4293
    #10;
    addra = 32'd137408;
    dina = {96'd0, 16'd51232, 16'd16111, 16'd45143, 16'd17486, 16'd53232, 16'd434, 16'd6874, 16'd65437, 16'd38902, 16'd33164}; // indx = 4294
    #10;
    addra = 32'd137440;
    dina = {96'd0, 16'd37937, 16'd56236, 16'd45223, 16'd25095, 16'd53172, 16'd21803, 16'd51769, 16'd32010, 16'd38165, 16'd59891}; // indx = 4295
    #10;
    addra = 32'd137472;
    dina = {96'd0, 16'd19223, 16'd48089, 16'd21356, 16'd41577, 16'd27693, 16'd4289, 16'd54124, 16'd4975, 16'd20598, 16'd848}; // indx = 4296
    #10;
    addra = 32'd137504;
    dina = {96'd0, 16'd53538, 16'd58302, 16'd44453, 16'd11190, 16'd35216, 16'd53785, 16'd45561, 16'd15887, 16'd64309, 16'd13160}; // indx = 4297
    #10;
    addra = 32'd137536;
    dina = {96'd0, 16'd45519, 16'd50943, 16'd10095, 16'd27729, 16'd57281, 16'd43488, 16'd52434, 16'd52552, 16'd902, 16'd58276}; // indx = 4298
    #10;
    addra = 32'd137568;
    dina = {96'd0, 16'd17517, 16'd8250, 16'd57173, 16'd16456, 16'd43718, 16'd30766, 16'd33862, 16'd42786, 16'd26875, 16'd23292}; // indx = 4299
    #10;
    addra = 32'd137600;
    dina = {96'd0, 16'd38260, 16'd24765, 16'd13221, 16'd44771, 16'd26576, 16'd8228, 16'd56823, 16'd46418, 16'd41616, 16'd12431}; // indx = 4300
    #10;
    addra = 32'd137632;
    dina = {96'd0, 16'd45170, 16'd50137, 16'd39131, 16'd12371, 16'd23159, 16'd56632, 16'd40501, 16'd23513, 16'd28170, 16'd54159}; // indx = 4301
    #10;
    addra = 32'd137664;
    dina = {96'd0, 16'd49791, 16'd30566, 16'd48094, 16'd42820, 16'd36269, 16'd23843, 16'd43255, 16'd42932, 16'd55824, 16'd24112}; // indx = 4302
    #10;
    addra = 32'd137696;
    dina = {96'd0, 16'd4902, 16'd11249, 16'd27092, 16'd53644, 16'd5539, 16'd16048, 16'd42188, 16'd32928, 16'd64629, 16'd65106}; // indx = 4303
    #10;
    addra = 32'd137728;
    dina = {96'd0, 16'd38779, 16'd50470, 16'd21187, 16'd4173, 16'd63764, 16'd60851, 16'd6411, 16'd41032, 16'd46921, 16'd54778}; // indx = 4304
    #10;
    addra = 32'd137760;
    dina = {96'd0, 16'd46293, 16'd36342, 16'd34635, 16'd13103, 16'd54983, 16'd36097, 16'd58521, 16'd20342, 16'd16689, 16'd65215}; // indx = 4305
    #10;
    addra = 32'd137792;
    dina = {96'd0, 16'd34917, 16'd51378, 16'd42678, 16'd64681, 16'd36104, 16'd46000, 16'd45108, 16'd42251, 16'd12850, 16'd52819}; // indx = 4306
    #10;
    addra = 32'd137824;
    dina = {96'd0, 16'd57658, 16'd21116, 16'd5831, 16'd43916, 16'd42593, 16'd60554, 16'd56959, 16'd43282, 16'd6971, 16'd26984}; // indx = 4307
    #10;
    addra = 32'd137856;
    dina = {96'd0, 16'd53224, 16'd50828, 16'd10031, 16'd1336, 16'd65130, 16'd5871, 16'd21679, 16'd62602, 16'd59386, 16'd11717}; // indx = 4308
    #10;
    addra = 32'd137888;
    dina = {96'd0, 16'd42717, 16'd8220, 16'd36164, 16'd15742, 16'd20725, 16'd7940, 16'd10382, 16'd49166, 16'd155, 16'd52126}; // indx = 4309
    #10;
    addra = 32'd137920;
    dina = {96'd0, 16'd58128, 16'd64108, 16'd9781, 16'd11860, 16'd1866, 16'd38561, 16'd12960, 16'd33454, 16'd3035, 16'd1481}; // indx = 4310
    #10;
    addra = 32'd137952;
    dina = {96'd0, 16'd53360, 16'd17894, 16'd1933, 16'd50451, 16'd23598, 16'd1183, 16'd48809, 16'd3592, 16'd48349, 16'd34803}; // indx = 4311
    #10;
    addra = 32'd137984;
    dina = {96'd0, 16'd7984, 16'd10274, 16'd45672, 16'd21394, 16'd6142, 16'd16592, 16'd32092, 16'd16323, 16'd46019, 16'd40356}; // indx = 4312
    #10;
    addra = 32'd138016;
    dina = {96'd0, 16'd17942, 16'd50463, 16'd55877, 16'd19981, 16'd58573, 16'd21373, 16'd17067, 16'd7733, 16'd58940, 16'd24836}; // indx = 4313
    #10;
    addra = 32'd138048;
    dina = {96'd0, 16'd20004, 16'd31138, 16'd47174, 16'd25622, 16'd15426, 16'd10591, 16'd26773, 16'd24409, 16'd8691, 16'd9298}; // indx = 4314
    #10;
    addra = 32'd138080;
    dina = {96'd0, 16'd7673, 16'd14334, 16'd20309, 16'd20229, 16'd21519, 16'd38550, 16'd32447, 16'd5528, 16'd34678, 16'd11028}; // indx = 4315
    #10;
    addra = 32'd138112;
    dina = {96'd0, 16'd42036, 16'd33367, 16'd59596, 16'd58563, 16'd39939, 16'd15757, 16'd31484, 16'd43367, 16'd21664, 16'd15919}; // indx = 4316
    #10;
    addra = 32'd138144;
    dina = {96'd0, 16'd37839, 16'd12467, 16'd11502, 16'd55233, 16'd33561, 16'd62538, 16'd24612, 16'd31482, 16'd47779, 16'd54176}; // indx = 4317
    #10;
    addra = 32'd138176;
    dina = {96'd0, 16'd42792, 16'd15187, 16'd19757, 16'd54812, 16'd51698, 16'd47542, 16'd61025, 16'd18373, 16'd4144, 16'd17752}; // indx = 4318
    #10;
    addra = 32'd138208;
    dina = {96'd0, 16'd50279, 16'd37599, 16'd20737, 16'd39907, 16'd23289, 16'd56078, 16'd52553, 16'd17482, 16'd4862, 16'd575}; // indx = 4319
    #10;
    addra = 32'd138240;
    dina = {96'd0, 16'd61349, 16'd20682, 16'd57883, 16'd6532, 16'd46170, 16'd58526, 16'd63344, 16'd29696, 16'd54939, 16'd8369}; // indx = 4320
    #10;
    addra = 32'd138272;
    dina = {96'd0, 16'd44470, 16'd54278, 16'd27296, 16'd32224, 16'd44812, 16'd29252, 16'd4228, 16'd18367, 16'd50427, 16'd18521}; // indx = 4321
    #10;
    addra = 32'd138304;
    dina = {96'd0, 16'd31734, 16'd29101, 16'd37295, 16'd64372, 16'd20231, 16'd4048, 16'd40161, 16'd42771, 16'd14725, 16'd21208}; // indx = 4322
    #10;
    addra = 32'd138336;
    dina = {96'd0, 16'd56705, 16'd2823, 16'd21179, 16'd19856, 16'd2905, 16'd61081, 16'd26637, 16'd12064, 16'd59213, 16'd64864}; // indx = 4323
    #10;
    addra = 32'd138368;
    dina = {96'd0, 16'd6352, 16'd5120, 16'd3148, 16'd36730, 16'd29818, 16'd41649, 16'd26868, 16'd49281, 16'd17489, 16'd42922}; // indx = 4324
    #10;
    addra = 32'd138400;
    dina = {96'd0, 16'd25923, 16'd23563, 16'd17084, 16'd26989, 16'd33369, 16'd18495, 16'd59150, 16'd12375, 16'd52903, 16'd63932}; // indx = 4325
    #10;
    addra = 32'd138432;
    dina = {96'd0, 16'd24391, 16'd7748, 16'd23901, 16'd6739, 16'd40762, 16'd25800, 16'd55271, 16'd2235, 16'd36568, 16'd22384}; // indx = 4326
    #10;
    addra = 32'd138464;
    dina = {96'd0, 16'd3923, 16'd65526, 16'd28245, 16'd20189, 16'd29107, 16'd62383, 16'd30467, 16'd57966, 16'd61079, 16'd30000}; // indx = 4327
    #10;
    addra = 32'd138496;
    dina = {96'd0, 16'd46195, 16'd36648, 16'd22280, 16'd671, 16'd17836, 16'd20870, 16'd19079, 16'd46152, 16'd60256, 16'd30015}; // indx = 4328
    #10;
    addra = 32'd138528;
    dina = {96'd0, 16'd30042, 16'd7552, 16'd59740, 16'd31576, 16'd62335, 16'd64685, 16'd48368, 16'd50966, 16'd46155, 16'd53043}; // indx = 4329
    #10;
    addra = 32'd138560;
    dina = {96'd0, 16'd49407, 16'd32654, 16'd65129, 16'd13770, 16'd30778, 16'd24424, 16'd27325, 16'd7146, 16'd47165, 16'd61164}; // indx = 4330
    #10;
    addra = 32'd138592;
    dina = {96'd0, 16'd8473, 16'd58178, 16'd15423, 16'd55426, 16'd51576, 16'd44705, 16'd42467, 16'd65385, 16'd41913, 16'd58106}; // indx = 4331
    #10;
    addra = 32'd138624;
    dina = {96'd0, 16'd24394, 16'd7111, 16'd42036, 16'd63744, 16'd32090, 16'd18491, 16'd26101, 16'd62631, 16'd20954, 16'd62854}; // indx = 4332
    #10;
    addra = 32'd138656;
    dina = {96'd0, 16'd4857, 16'd23750, 16'd51432, 16'd23785, 16'd18570, 16'd51031, 16'd51343, 16'd60127, 16'd54824, 16'd20138}; // indx = 4333
    #10;
    addra = 32'd138688;
    dina = {96'd0, 16'd40129, 16'd51856, 16'd25602, 16'd43201, 16'd54415, 16'd53888, 16'd44673, 16'd1445, 16'd18010, 16'd26113}; // indx = 4334
    #10;
    addra = 32'd138720;
    dina = {96'd0, 16'd3032, 16'd40483, 16'd35864, 16'd18549, 16'd28178, 16'd58199, 16'd59267, 16'd64027, 16'd44481, 16'd59545}; // indx = 4335
    #10;
    addra = 32'd138752;
    dina = {96'd0, 16'd1339, 16'd16414, 16'd35418, 16'd45723, 16'd10185, 16'd56498, 16'd64466, 16'd33536, 16'd4114, 16'd6533}; // indx = 4336
    #10;
    addra = 32'd138784;
    dina = {96'd0, 16'd17675, 16'd14256, 16'd59139, 16'd19337, 16'd30282, 16'd9734, 16'd34123, 16'd43127, 16'd56501, 16'd28798}; // indx = 4337
    #10;
    addra = 32'd138816;
    dina = {96'd0, 16'd58670, 16'd20425, 16'd57628, 16'd38856, 16'd3376, 16'd53543, 16'd63224, 16'd37295, 16'd50969, 16'd29572}; // indx = 4338
    #10;
    addra = 32'd138848;
    dina = {96'd0, 16'd39478, 16'd42617, 16'd31024, 16'd32540, 16'd15748, 16'd8055, 16'd29017, 16'd61499, 16'd24280, 16'd33460}; // indx = 4339
    #10;
    addra = 32'd138880;
    dina = {96'd0, 16'd54301, 16'd23193, 16'd54571, 16'd27924, 16'd25106, 16'd24870, 16'd21092, 16'd35719, 16'd44094, 16'd49526}; // indx = 4340
    #10;
    addra = 32'd138912;
    dina = {96'd0, 16'd43001, 16'd23517, 16'd50504, 16'd45952, 16'd35082, 16'd27575, 16'd24251, 16'd51600, 16'd61530, 16'd26487}; // indx = 4341
    #10;
    addra = 32'd138944;
    dina = {96'd0, 16'd51695, 16'd65389, 16'd6442, 16'd17469, 16'd68, 16'd65445, 16'd43451, 16'd51911, 16'd41030, 16'd1146}; // indx = 4342
    #10;
    addra = 32'd138976;
    dina = {96'd0, 16'd33644, 16'd2996, 16'd37814, 16'd41967, 16'd49533, 16'd45684, 16'd41328, 16'd58177, 16'd58123, 16'd57274}; // indx = 4343
    #10;
    addra = 32'd139008;
    dina = {96'd0, 16'd3023, 16'd12647, 16'd62514, 16'd7008, 16'd54440, 16'd60013, 16'd1565, 16'd60420, 16'd39667, 16'd25498}; // indx = 4344
    #10;
    addra = 32'd139040;
    dina = {96'd0, 16'd20, 16'd36759, 16'd50078, 16'd64734, 16'd24259, 16'd16153, 16'd47026, 16'd56311, 16'd3742, 16'd49535}; // indx = 4345
    #10;
    addra = 32'd139072;
    dina = {96'd0, 16'd26722, 16'd22933, 16'd817, 16'd124, 16'd4249, 16'd52486, 16'd33759, 16'd4117, 16'd19702, 16'd31250}; // indx = 4346
    #10;
    addra = 32'd139104;
    dina = {96'd0, 16'd60014, 16'd60983, 16'd64803, 16'd22483, 16'd65508, 16'd12987, 16'd37020, 16'd23110, 16'd6095, 16'd18060}; // indx = 4347
    #10;
    addra = 32'd139136;
    dina = {96'd0, 16'd22646, 16'd12478, 16'd22357, 16'd21529, 16'd41546, 16'd61346, 16'd19152, 16'd8029, 16'd43463, 16'd3549}; // indx = 4348
    #10;
    addra = 32'd139168;
    dina = {96'd0, 16'd17365, 16'd6571, 16'd3492, 16'd56370, 16'd65474, 16'd28528, 16'd49361, 16'd23924, 16'd39935, 16'd2489}; // indx = 4349
    #10;
    addra = 32'd139200;
    dina = {96'd0, 16'd9839, 16'd881, 16'd5037, 16'd24470, 16'd47801, 16'd21307, 16'd14647, 16'd12313, 16'd53218, 16'd59363}; // indx = 4350
    #10;
    addra = 32'd139232;
    dina = {96'd0, 16'd35694, 16'd39814, 16'd58987, 16'd25557, 16'd34532, 16'd65153, 16'd18406, 16'd31205, 16'd55094, 16'd3000}; // indx = 4351
    #10;
    addra = 32'd139264;
    dina = {96'd0, 16'd53218, 16'd48829, 16'd55082, 16'd1391, 16'd39041, 16'd3560, 16'd42412, 16'd10499, 16'd40997, 16'd33084}; // indx = 4352
    #10;
    addra = 32'd139296;
    dina = {96'd0, 16'd8968, 16'd49969, 16'd60485, 16'd27946, 16'd63697, 16'd46009, 16'd51606, 16'd8120, 16'd45981, 16'd37043}; // indx = 4353
    #10;
    addra = 32'd139328;
    dina = {96'd0, 16'd7671, 16'd43084, 16'd42137, 16'd28848, 16'd33880, 16'd31905, 16'd44869, 16'd48653, 16'd43830, 16'd6464}; // indx = 4354
    #10;
    addra = 32'd139360;
    dina = {96'd0, 16'd13147, 16'd36826, 16'd21501, 16'd19924, 16'd38278, 16'd7865, 16'd64921, 16'd2639, 16'd59477, 16'd57821}; // indx = 4355
    #10;
    addra = 32'd139392;
    dina = {96'd0, 16'd4251, 16'd46288, 16'd32776, 16'd52288, 16'd50723, 16'd24502, 16'd33824, 16'd43336, 16'd39862, 16'd39257}; // indx = 4356
    #10;
    addra = 32'd139424;
    dina = {96'd0, 16'd25643, 16'd9352, 16'd8975, 16'd712, 16'd11880, 16'd34510, 16'd40426, 16'd35235, 16'd60449, 16'd11171}; // indx = 4357
    #10;
    addra = 32'd139456;
    dina = {96'd0, 16'd37633, 16'd59860, 16'd9407, 16'd30966, 16'd63473, 16'd2054, 16'd11350, 16'd17250, 16'd46154, 16'd2924}; // indx = 4358
    #10;
    addra = 32'd139488;
    dina = {96'd0, 16'd10319, 16'd41102, 16'd35855, 16'd9424, 16'd31164, 16'd46920, 16'd35368, 16'd59303, 16'd18975, 16'd55}; // indx = 4359
    #10;
    addra = 32'd139520;
    dina = {96'd0, 16'd39280, 16'd58309, 16'd52346, 16'd22260, 16'd12656, 16'd37225, 16'd35665, 16'd21719, 16'd11575, 16'd30904}; // indx = 4360
    #10;
    addra = 32'd139552;
    dina = {96'd0, 16'd44511, 16'd7532, 16'd61428, 16'd28662, 16'd2629, 16'd40278, 16'd26039, 16'd44510, 16'd26923, 16'd2637}; // indx = 4361
    #10;
    addra = 32'd139584;
    dina = {96'd0, 16'd21265, 16'd46465, 16'd13021, 16'd49874, 16'd18502, 16'd21738, 16'd57126, 16'd49230, 16'd15823, 16'd16642}; // indx = 4362
    #10;
    addra = 32'd139616;
    dina = {96'd0, 16'd52724, 16'd54409, 16'd53251, 16'd24154, 16'd54299, 16'd61759, 16'd61599, 16'd51918, 16'd58402, 16'd3266}; // indx = 4363
    #10;
    addra = 32'd139648;
    dina = {96'd0, 16'd13925, 16'd5615, 16'd2087, 16'd49984, 16'd20054, 16'd24760, 16'd55923, 16'd686, 16'd7842, 16'd31766}; // indx = 4364
    #10;
    addra = 32'd139680;
    dina = {96'd0, 16'd35872, 16'd11009, 16'd10296, 16'd965, 16'd43925, 16'd32698, 16'd258, 16'd24157, 16'd24309, 16'd53355}; // indx = 4365
    #10;
    addra = 32'd139712;
    dina = {96'd0, 16'd11264, 16'd37592, 16'd23699, 16'd35318, 16'd53622, 16'd46546, 16'd26548, 16'd7329, 16'd60281, 16'd25998}; // indx = 4366
    #10;
    addra = 32'd139744;
    dina = {96'd0, 16'd65221, 16'd37199, 16'd62876, 16'd36943, 16'd38763, 16'd8696, 16'd20893, 16'd26728, 16'd7411, 16'd30916}; // indx = 4367
    #10;
    addra = 32'd139776;
    dina = {96'd0, 16'd57937, 16'd9081, 16'd24678, 16'd56667, 16'd16999, 16'd16093, 16'd10995, 16'd7127, 16'd40613, 16'd10738}; // indx = 4368
    #10;
    addra = 32'd139808;
    dina = {96'd0, 16'd37624, 16'd863, 16'd60216, 16'd39556, 16'd44792, 16'd24506, 16'd35263, 16'd37374, 16'd8405, 16'd1289}; // indx = 4369
    #10;
    addra = 32'd139840;
    dina = {96'd0, 16'd17573, 16'd11143, 16'd22901, 16'd27624, 16'd25239, 16'd65275, 16'd65129, 16'd20284, 16'd24361, 16'd12555}; // indx = 4370
    #10;
    addra = 32'd139872;
    dina = {96'd0, 16'd42993, 16'd55822, 16'd29680, 16'd22808, 16'd50098, 16'd21379, 16'd20455, 16'd2880, 16'd18843, 16'd35667}; // indx = 4371
    #10;
    addra = 32'd139904;
    dina = {96'd0, 16'd10837, 16'd4433, 16'd27733, 16'd31966, 16'd616, 16'd25089, 16'd55143, 16'd4252, 16'd4157, 16'd35997}; // indx = 4372
    #10;
    addra = 32'd139936;
    dina = {96'd0, 16'd14768, 16'd52403, 16'd16082, 16'd52339, 16'd20180, 16'd42395, 16'd9519, 16'd18149, 16'd55501, 16'd8702}; // indx = 4373
    #10;
    addra = 32'd139968;
    dina = {96'd0, 16'd4125, 16'd17926, 16'd7323, 16'd48387, 16'd40177, 16'd36518, 16'd54552, 16'd14043, 16'd54335, 16'd9912}; // indx = 4374
    #10;
    addra = 32'd140000;
    dina = {96'd0, 16'd48614, 16'd47487, 16'd34456, 16'd31368, 16'd41440, 16'd60512, 16'd19890, 16'd42227, 16'd16950, 16'd16774}; // indx = 4375
    #10;
    addra = 32'd140032;
    dina = {96'd0, 16'd20741, 16'd29246, 16'd53596, 16'd58178, 16'd12181, 16'd43490, 16'd32147, 16'd38324, 16'd57481, 16'd36257}; // indx = 4376
    #10;
    addra = 32'd140064;
    dina = {96'd0, 16'd33511, 16'd24441, 16'd23089, 16'd59096, 16'd931, 16'd30125, 16'd29628, 16'd65267, 16'd18185, 16'd18282}; // indx = 4377
    #10;
    addra = 32'd140096;
    dina = {96'd0, 16'd5766, 16'd34181, 16'd42803, 16'd14097, 16'd6383, 16'd52608, 16'd35508, 16'd64381, 16'd59416, 16'd35738}; // indx = 4378
    #10;
    addra = 32'd140128;
    dina = {96'd0, 16'd14483, 16'd54899, 16'd36234, 16'd57025, 16'd30113, 16'd52928, 16'd37956, 16'd25417, 16'd63737, 16'd15020}; // indx = 4379
    #10;
    addra = 32'd140160;
    dina = {96'd0, 16'd13411, 16'd54358, 16'd30503, 16'd12709, 16'd65069, 16'd40533, 16'd23488, 16'd63163, 16'd48062, 16'd26158}; // indx = 4380
    #10;
    addra = 32'd140192;
    dina = {96'd0, 16'd1443, 16'd51978, 16'd19429, 16'd7426, 16'd3160, 16'd39052, 16'd38297, 16'd63817, 16'd17747, 16'd32097}; // indx = 4381
    #10;
    addra = 32'd140224;
    dina = {96'd0, 16'd4875, 16'd30150, 16'd34441, 16'd59346, 16'd19469, 16'd29425, 16'd5431, 16'd29773, 16'd51197, 16'd26191}; // indx = 4382
    #10;
    addra = 32'd140256;
    dina = {96'd0, 16'd686, 16'd45574, 16'd45057, 16'd10668, 16'd21767, 16'd58207, 16'd55987, 16'd10478, 16'd37997, 16'd48469}; // indx = 4383
    #10;
    addra = 32'd140288;
    dina = {96'd0, 16'd5834, 16'd59363, 16'd59441, 16'd21249, 16'd18803, 16'd32621, 16'd45732, 16'd40448, 16'd45224, 16'd48628}; // indx = 4384
    #10;
    addra = 32'd140320;
    dina = {96'd0, 16'd46691, 16'd26054, 16'd13729, 16'd61421, 16'd1396, 16'd43561, 16'd30693, 16'd51736, 16'd6834, 16'd60675}; // indx = 4385
    #10;
    addra = 32'd140352;
    dina = {96'd0, 16'd26063, 16'd37751, 16'd43866, 16'd27890, 16'd16436, 16'd54778, 16'd26972, 16'd40050, 16'd19282, 16'd44500}; // indx = 4386
    #10;
    addra = 32'd140384;
    dina = {96'd0, 16'd22749, 16'd38941, 16'd6640, 16'd9692, 16'd34113, 16'd28989, 16'd34265, 16'd53344, 16'd31031, 16'd63181}; // indx = 4387
    #10;
    addra = 32'd140416;
    dina = {96'd0, 16'd12186, 16'd62801, 16'd55990, 16'd60798, 16'd63829, 16'd54935, 16'd38555, 16'd52724, 16'd10436, 16'd11252}; // indx = 4388
    #10;
    addra = 32'd140448;
    dina = {96'd0, 16'd16818, 16'd11781, 16'd18112, 16'd19039, 16'd64740, 16'd55741, 16'd14068, 16'd1737, 16'd61615, 16'd23884}; // indx = 4389
    #10;
    addra = 32'd140480;
    dina = {96'd0, 16'd13775, 16'd48396, 16'd61288, 16'd4244, 16'd41367, 16'd5460, 16'd54694, 16'd51224, 16'd10788, 16'd62213}; // indx = 4390
    #10;
    addra = 32'd140512;
    dina = {96'd0, 16'd10051, 16'd8206, 16'd18486, 16'd36740, 16'd9764, 16'd23871, 16'd31911, 16'd60113, 16'd22974, 16'd34108}; // indx = 4391
    #10;
    addra = 32'd140544;
    dina = {96'd0, 16'd48507, 16'd53195, 16'd46479, 16'd20296, 16'd10592, 16'd14103, 16'd37329, 16'd26678, 16'd59157, 16'd28872}; // indx = 4392
    #10;
    addra = 32'd140576;
    dina = {96'd0, 16'd49747, 16'd40083, 16'd63202, 16'd22651, 16'd28323, 16'd30207, 16'd4456, 16'd16801, 16'd50425, 16'd8644}; // indx = 4393
    #10;
    addra = 32'd140608;
    dina = {96'd0, 16'd45438, 16'd65144, 16'd12704, 16'd62617, 16'd54261, 16'd37528, 16'd57691, 16'd59961, 16'd59484, 16'd43719}; // indx = 4394
    #10;
    addra = 32'd140640;
    dina = {96'd0, 16'd46239, 16'd4359, 16'd1749, 16'd35909, 16'd33562, 16'd50931, 16'd43554, 16'd29447, 16'd2127, 16'd25821}; // indx = 4395
    #10;
    addra = 32'd140672;
    dina = {96'd0, 16'd19195, 16'd31511, 16'd26080, 16'd44664, 16'd40380, 16'd32283, 16'd17028, 16'd35044, 16'd52714, 16'd47348}; // indx = 4396
    #10;
    addra = 32'd140704;
    dina = {96'd0, 16'd6513, 16'd30685, 16'd36432, 16'd12716, 16'd8083, 16'd2783, 16'd22853, 16'd30934, 16'd35708, 16'd58463}; // indx = 4397
    #10;
    addra = 32'd140736;
    dina = {96'd0, 16'd27272, 16'd58497, 16'd5957, 16'd38378, 16'd11578, 16'd21420, 16'd32782, 16'd15030, 16'd33310, 16'd40661}; // indx = 4398
    #10;
    addra = 32'd140768;
    dina = {96'd0, 16'd9234, 16'd30579, 16'd63258, 16'd46526, 16'd10283, 16'd51615, 16'd10458, 16'd19464, 16'd27629, 16'd7236}; // indx = 4399
    #10;
    addra = 32'd140800;
    dina = {96'd0, 16'd33949, 16'd5787, 16'd40707, 16'd47492, 16'd39179, 16'd26151, 16'd18196, 16'd37383, 16'd15847, 16'd132}; // indx = 4400
    #10;
    addra = 32'd140832;
    dina = {96'd0, 16'd12483, 16'd1223, 16'd23091, 16'd2227, 16'd12019, 16'd51198, 16'd26200, 16'd24690, 16'd519, 16'd25398}; // indx = 4401
    #10;
    addra = 32'd140864;
    dina = {96'd0, 16'd44368, 16'd41726, 16'd47616, 16'd33521, 16'd61705, 16'd11239, 16'd44397, 16'd24716, 16'd63445, 16'd60560}; // indx = 4402
    #10;
    addra = 32'd140896;
    dina = {96'd0, 16'd50719, 16'd8955, 16'd40057, 16'd49185, 16'd28751, 16'd8889, 16'd47872, 16'd48232, 16'd38884, 16'd33608}; // indx = 4403
    #10;
    addra = 32'd140928;
    dina = {96'd0, 16'd26017, 16'd1236, 16'd30717, 16'd3034, 16'd54217, 16'd12043, 16'd47946, 16'd15031, 16'd28234, 16'd9161}; // indx = 4404
    #10;
    addra = 32'd140960;
    dina = {96'd0, 16'd52123, 16'd3016, 16'd47589, 16'd16266, 16'd28878, 16'd31990, 16'd61764, 16'd43558, 16'd1891, 16'd31483}; // indx = 4405
    #10;
    addra = 32'd140992;
    dina = {96'd0, 16'd51812, 16'd18702, 16'd59976, 16'd31481, 16'd22928, 16'd14698, 16'd31495, 16'd62206, 16'd48072, 16'd6669}; // indx = 4406
    #10;
    addra = 32'd141024;
    dina = {96'd0, 16'd35435, 16'd31814, 16'd34274, 16'd53614, 16'd29356, 16'd59903, 16'd41523, 16'd18808, 16'd13398, 16'd6030}; // indx = 4407
    #10;
    addra = 32'd141056;
    dina = {96'd0, 16'd49511, 16'd17863, 16'd46421, 16'd462, 16'd23718, 16'd11379, 16'd55590, 16'd44408, 16'd9868, 16'd62051}; // indx = 4408
    #10;
    addra = 32'd141088;
    dina = {96'd0, 16'd53318, 16'd20586, 16'd7727, 16'd21334, 16'd30595, 16'd22736, 16'd60573, 16'd61813, 16'd27084, 16'd55415}; // indx = 4409
    #10;
    addra = 32'd141120;
    dina = {96'd0, 16'd47046, 16'd17932, 16'd45028, 16'd45586, 16'd5473, 16'd40055, 16'd32393, 16'd55466, 16'd1622, 16'd12991}; // indx = 4410
    #10;
    addra = 32'd141152;
    dina = {96'd0, 16'd6729, 16'd65353, 16'd13167, 16'd50005, 16'd60387, 16'd21295, 16'd26054, 16'd22335, 16'd44914, 16'd31696}; // indx = 4411
    #10;
    addra = 32'd141184;
    dina = {96'd0, 16'd29293, 16'd11218, 16'd65346, 16'd43772, 16'd48934, 16'd21080, 16'd39273, 16'd21923, 16'd42842, 16'd44301}; // indx = 4412
    #10;
    addra = 32'd141216;
    dina = {96'd0, 16'd62339, 16'd47660, 16'd23882, 16'd17211, 16'd24299, 16'd10903, 16'd35235, 16'd56537, 16'd56338, 16'd5407}; // indx = 4413
    #10;
    addra = 32'd141248;
    dina = {96'd0, 16'd28853, 16'd44913, 16'd58559, 16'd40334, 16'd10546, 16'd38305, 16'd22679, 16'd1240, 16'd53692, 16'd13178}; // indx = 4414
    #10;
    addra = 32'd141280;
    dina = {96'd0, 16'd13066, 16'd28141, 16'd55283, 16'd3183, 16'd60854, 16'd42589, 16'd59090, 16'd43655, 16'd52576, 16'd39957}; // indx = 4415
    #10;
    addra = 32'd141312;
    dina = {96'd0, 16'd58256, 16'd52150, 16'd20561, 16'd21592, 16'd43252, 16'd1667, 16'd10282, 16'd28129, 16'd10275, 16'd14353}; // indx = 4416
    #10;
    addra = 32'd141344;
    dina = {96'd0, 16'd3624, 16'd49598, 16'd88, 16'd39856, 16'd53553, 16'd64853, 16'd63506, 16'd37938, 16'd35404, 16'd4465}; // indx = 4417
    #10;
    addra = 32'd141376;
    dina = {96'd0, 16'd51685, 16'd8594, 16'd7436, 16'd45579, 16'd11441, 16'd47983, 16'd41684, 16'd47867, 16'd50966, 16'd37580}; // indx = 4418
    #10;
    addra = 32'd141408;
    dina = {96'd0, 16'd37414, 16'd55723, 16'd671, 16'd19939, 16'd22339, 16'd2515, 16'd3418, 16'd49534, 16'd4652, 16'd64125}; // indx = 4419
    #10;
    addra = 32'd141440;
    dina = {96'd0, 16'd46572, 16'd19468, 16'd58079, 16'd16441, 16'd29167, 16'd29963, 16'd61319, 16'd80, 16'd54386, 16'd51911}; // indx = 4420
    #10;
    addra = 32'd141472;
    dina = {96'd0, 16'd47591, 16'd4647, 16'd33447, 16'd31304, 16'd19509, 16'd36583, 16'd31331, 16'd41015, 16'd13407, 16'd1770}; // indx = 4421
    #10;
    addra = 32'd141504;
    dina = {96'd0, 16'd23686, 16'd54517, 16'd24882, 16'd41991, 16'd11946, 16'd880, 16'd44325, 16'd18903, 16'd2357, 16'd56988}; // indx = 4422
    #10;
    addra = 32'd141536;
    dina = {96'd0, 16'd57058, 16'd57634, 16'd16779, 16'd26915, 16'd64228, 16'd56842, 16'd55131, 16'd21283, 16'd35788, 16'd62963}; // indx = 4423
    #10;
    addra = 32'd141568;
    dina = {96'd0, 16'd38545, 16'd9615, 16'd19770, 16'd25186, 16'd58034, 16'd25760, 16'd36019, 16'd57082, 16'd36056, 16'd56852}; // indx = 4424
    #10;
    addra = 32'd141600;
    dina = {96'd0, 16'd34603, 16'd14913, 16'd32571, 16'd35234, 16'd34233, 16'd31983, 16'd63087, 16'd43332, 16'd33555, 16'd8282}; // indx = 4425
    #10;
    addra = 32'd141632;
    dina = {96'd0, 16'd22310, 16'd55015, 16'd2469, 16'd10819, 16'd34482, 16'd44335, 16'd51054, 16'd7150, 16'd41603, 16'd25576}; // indx = 4426
    #10;
    addra = 32'd141664;
    dina = {96'd0, 16'd50018, 16'd60144, 16'd9461, 16'd41168, 16'd22094, 16'd20744, 16'd29288, 16'd46932, 16'd2267, 16'd15591}; // indx = 4427
    #10;
    addra = 32'd141696;
    dina = {96'd0, 16'd2166, 16'd25231, 16'd18499, 16'd42942, 16'd22521, 16'd27401, 16'd61667, 16'd14518, 16'd63615, 16'd45718}; // indx = 4428
    #10;
    addra = 32'd141728;
    dina = {96'd0, 16'd17052, 16'd5520, 16'd48578, 16'd19099, 16'd33228, 16'd57184, 16'd63238, 16'd37057, 16'd10878, 16'd24955}; // indx = 4429
    #10;
    addra = 32'd141760;
    dina = {96'd0, 16'd46716, 16'd47515, 16'd30447, 16'd19610, 16'd29666, 16'd26011, 16'd14066, 16'd18331, 16'd55882, 16'd57205}; // indx = 4430
    #10;
    addra = 32'd141792;
    dina = {96'd0, 16'd43763, 16'd39681, 16'd60178, 16'd54514, 16'd51605, 16'd10391, 16'd59631, 16'd16722, 16'd10059, 16'd28266}; // indx = 4431
    #10;
    addra = 32'd141824;
    dina = {96'd0, 16'd19435, 16'd62622, 16'd23553, 16'd22760, 16'd1258, 16'd11762, 16'd55581, 16'd55072, 16'd20007, 16'd4542}; // indx = 4432
    #10;
    addra = 32'd141856;
    dina = {96'd0, 16'd52002, 16'd64888, 16'd35254, 16'd38096, 16'd18855, 16'd31205, 16'd50257, 16'd36965, 16'd53512, 16'd14572}; // indx = 4433
    #10;
    addra = 32'd141888;
    dina = {96'd0, 16'd45666, 16'd52118, 16'd55297, 16'd339, 16'd13127, 16'd17724, 16'd31775, 16'd10349, 16'd47843, 16'd26642}; // indx = 4434
    #10;
    addra = 32'd141920;
    dina = {96'd0, 16'd24785, 16'd40103, 16'd21655, 16'd57105, 16'd2393, 16'd35600, 16'd41301, 16'd60806, 16'd61903, 16'd22442}; // indx = 4435
    #10;
    addra = 32'd141952;
    dina = {96'd0, 16'd40202, 16'd1678, 16'd21525, 16'd2148, 16'd2813, 16'd47503, 16'd24471, 16'd23043, 16'd28366, 16'd43148}; // indx = 4436
    #10;
    addra = 32'd141984;
    dina = {96'd0, 16'd39648, 16'd43166, 16'd15087, 16'd56092, 16'd24658, 16'd43654, 16'd47891, 16'd60863, 16'd64344, 16'd2832}; // indx = 4437
    #10;
    addra = 32'd142016;
    dina = {96'd0, 16'd11983, 16'd268, 16'd1401, 16'd48413, 16'd47922, 16'd28832, 16'd51125, 16'd57774, 16'd21197, 16'd64369}; // indx = 4438
    #10;
    addra = 32'd142048;
    dina = {96'd0, 16'd46057, 16'd20781, 16'd36650, 16'd55909, 16'd13290, 16'd460, 16'd47493, 16'd12062, 16'd11436, 16'd4400}; // indx = 4439
    #10;
    addra = 32'd142080;
    dina = {96'd0, 16'd17158, 16'd15374, 16'd51360, 16'd9791, 16'd39359, 16'd59013, 16'd25172, 16'd40848, 16'd40219, 16'd53558}; // indx = 4440
    #10;
    addra = 32'd142112;
    dina = {96'd0, 16'd32913, 16'd59820, 16'd2774, 16'd19324, 16'd24580, 16'd26363, 16'd50094, 16'd48599, 16'd51218, 16'd36078}; // indx = 4441
    #10;
    addra = 32'd142144;
    dina = {96'd0, 16'd59142, 16'd26046, 16'd53288, 16'd50996, 16'd53768, 16'd59802, 16'd7905, 16'd21819, 16'd51266, 16'd44201}; // indx = 4442
    #10;
    addra = 32'd142176;
    dina = {96'd0, 16'd42820, 16'd54424, 16'd65450, 16'd57573, 16'd58249, 16'd34867, 16'd65278, 16'd14465, 16'd61673, 16'd12677}; // indx = 4443
    #10;
    addra = 32'd142208;
    dina = {96'd0, 16'd1499, 16'd59621, 16'd46651, 16'd2426, 16'd62851, 16'd6777, 16'd52742, 16'd12303, 16'd34564, 16'd25548}; // indx = 4444
    #10;
    addra = 32'd142240;
    dina = {96'd0, 16'd54916, 16'd41613, 16'd9996, 16'd8349, 16'd49880, 16'd14051, 16'd4908, 16'd5254, 16'd56187, 16'd40843}; // indx = 4445
    #10;
    addra = 32'd142272;
    dina = {96'd0, 16'd57001, 16'd51797, 16'd32753, 16'd16734, 16'd10593, 16'd52103, 16'd13021, 16'd53467, 16'd30070, 16'd4619}; // indx = 4446
    #10;
    addra = 32'd142304;
    dina = {96'd0, 16'd5868, 16'd50848, 16'd9760, 16'd11378, 16'd31264, 16'd10513, 16'd7353, 16'd23825, 16'd48489, 16'd37982}; // indx = 4447
    #10;
    addra = 32'd142336;
    dina = {96'd0, 16'd10973, 16'd34556, 16'd60892, 16'd35475, 16'd61747, 16'd20755, 16'd11327, 16'd24810, 16'd61643, 16'd23294}; // indx = 4448
    #10;
    addra = 32'd142368;
    dina = {96'd0, 16'd7639, 16'd30311, 16'd31759, 16'd7502, 16'd21215, 16'd32973, 16'd65260, 16'd20746, 16'd61274, 16'd24770}; // indx = 4449
    #10;
    addra = 32'd142400;
    dina = {96'd0, 16'd25491, 16'd58905, 16'd55741, 16'd7678, 16'd38870, 16'd44870, 16'd25698, 16'd39695, 16'd27755, 16'd38370}; // indx = 4450
    #10;
    addra = 32'd142432;
    dina = {96'd0, 16'd61795, 16'd1033, 16'd45095, 16'd58539, 16'd14240, 16'd14589, 16'd8442, 16'd3718, 16'd45550, 16'd23804}; // indx = 4451
    #10;
    addra = 32'd142464;
    dina = {96'd0, 16'd19028, 16'd925, 16'd53960, 16'd62952, 16'd35856, 16'd3697, 16'd34139, 16'd13140, 16'd37557, 16'd14383}; // indx = 4452
    #10;
    addra = 32'd142496;
    dina = {96'd0, 16'd53986, 16'd64848, 16'd52531, 16'd62712, 16'd27247, 16'd34276, 16'd62765, 16'd3663, 16'd20609, 16'd29117}; // indx = 4453
    #10;
    addra = 32'd142528;
    dina = {96'd0, 16'd62090, 16'd22128, 16'd7398, 16'd20249, 16'd60408, 16'd60009, 16'd61602, 16'd39779, 16'd58918, 16'd60159}; // indx = 4454
    #10;
    addra = 32'd142560;
    dina = {96'd0, 16'd33598, 16'd16149, 16'd26357, 16'd59522, 16'd11524, 16'd4736, 16'd28875, 16'd268, 16'd47308, 16'd40492}; // indx = 4455
    #10;
    addra = 32'd142592;
    dina = {96'd0, 16'd22109, 16'd25259, 16'd21180, 16'd10978, 16'd4640, 16'd22040, 16'd45460, 16'd25442, 16'd46065, 16'd2577}; // indx = 4456
    #10;
    addra = 32'd142624;
    dina = {96'd0, 16'd60340, 16'd49527, 16'd47220, 16'd44952, 16'd29255, 16'd49715, 16'd22370, 16'd63620, 16'd53565, 16'd30244}; // indx = 4457
    #10;
    addra = 32'd142656;
    dina = {96'd0, 16'd34786, 16'd13287, 16'd27752, 16'd16358, 16'd44494, 16'd356, 16'd38156, 16'd8846, 16'd28322, 16'd41406}; // indx = 4458
    #10;
    addra = 32'd142688;
    dina = {96'd0, 16'd3482, 16'd57426, 16'd61452, 16'd42778, 16'd38285, 16'd26676, 16'd5506, 16'd9515, 16'd34811, 16'd3559}; // indx = 4459
    #10;
    addra = 32'd142720;
    dina = {96'd0, 16'd8030, 16'd45718, 16'd3509, 16'd33708, 16'd18632, 16'd8916, 16'd61783, 16'd34830, 16'd21640, 16'd56212}; // indx = 4460
    #10;
    addra = 32'd142752;
    dina = {96'd0, 16'd53557, 16'd59114, 16'd62362, 16'd4939, 16'd64804, 16'd55923, 16'd64889, 16'd16093, 16'd6325, 16'd28144}; // indx = 4461
    #10;
    addra = 32'd142784;
    dina = {96'd0, 16'd20584, 16'd4951, 16'd19755, 16'd56001, 16'd49996, 16'd8334, 16'd45379, 16'd43057, 16'd39379, 16'd11072}; // indx = 4462
    #10;
    addra = 32'd142816;
    dina = {96'd0, 16'd24030, 16'd53570, 16'd2007, 16'd19188, 16'd2335, 16'd9030, 16'd5153, 16'd22272, 16'd10382, 16'd64219}; // indx = 4463
    #10;
    addra = 32'd142848;
    dina = {96'd0, 16'd14567, 16'd20269, 16'd5497, 16'd45505, 16'd189, 16'd59867, 16'd21285, 16'd32022, 16'd29673, 16'd5873}; // indx = 4464
    #10;
    addra = 32'd142880;
    dina = {96'd0, 16'd8320, 16'd2189, 16'd28663, 16'd54922, 16'd31794, 16'd30743, 16'd8967, 16'd28084, 16'd26886, 16'd61818}; // indx = 4465
    #10;
    addra = 32'd142912;
    dina = {96'd0, 16'd17314, 16'd31659, 16'd21305, 16'd60565, 16'd7462, 16'd23421, 16'd13364, 16'd47579, 16'd58496, 16'd31921}; // indx = 4466
    #10;
    addra = 32'd142944;
    dina = {96'd0, 16'd49644, 16'd6084, 16'd61544, 16'd10916, 16'd656, 16'd46351, 16'd42732, 16'd10434, 16'd45682, 16'd46542}; // indx = 4467
    #10;
    addra = 32'd142976;
    dina = {96'd0, 16'd48629, 16'd29609, 16'd64725, 16'd23936, 16'd44150, 16'd31228, 16'd56314, 16'd21278, 16'd59746, 16'd25501}; // indx = 4468
    #10;
    addra = 32'd143008;
    dina = {96'd0, 16'd49704, 16'd12975, 16'd42209, 16'd34213, 16'd33709, 16'd64250, 16'd35726, 16'd62213, 16'd100, 16'd15550}; // indx = 4469
    #10;
    addra = 32'd143040;
    dina = {96'd0, 16'd37287, 16'd2900, 16'd45031, 16'd34384, 16'd34827, 16'd28045, 16'd41187, 16'd2430, 16'd46521, 16'd21951}; // indx = 4470
    #10;
    addra = 32'd143072;
    dina = {96'd0, 16'd2115, 16'd47600, 16'd62050, 16'd934, 16'd46689, 16'd43832, 16'd1322, 16'd33186, 16'd11181, 16'd3517}; // indx = 4471
    #10;
    addra = 32'd143104;
    dina = {96'd0, 16'd8615, 16'd34804, 16'd63717, 16'd3554, 16'd50494, 16'd33600, 16'd49927, 16'd12830, 16'd34572, 16'd2774}; // indx = 4472
    #10;
    addra = 32'd143136;
    dina = {96'd0, 16'd30408, 16'd49253, 16'd19289, 16'd46694, 16'd38655, 16'd42816, 16'd56569, 16'd326, 16'd36428, 16'd38184}; // indx = 4473
    #10;
    addra = 32'd143168;
    dina = {96'd0, 16'd51311, 16'd25945, 16'd44087, 16'd25053, 16'd44946, 16'd12233, 16'd19675, 16'd28635, 16'd52752, 16'd55304}; // indx = 4474
    #10;
    addra = 32'd143200;
    dina = {96'd0, 16'd26935, 16'd18220, 16'd16532, 16'd54230, 16'd19009, 16'd27067, 16'd54438, 16'd13815, 16'd18954, 16'd38362}; // indx = 4475
    #10;
    addra = 32'd143232;
    dina = {96'd0, 16'd14364, 16'd26779, 16'd7428, 16'd4566, 16'd38848, 16'd13818, 16'd6224, 16'd44616, 16'd6074, 16'd10824}; // indx = 4476
    #10;
    addra = 32'd143264;
    dina = {96'd0, 16'd51467, 16'd53976, 16'd27748, 16'd47571, 16'd3575, 16'd28830, 16'd46077, 16'd19697, 16'd39784, 16'd22773}; // indx = 4477
    #10;
    addra = 32'd143296;
    dina = {96'd0, 16'd14317, 16'd45188, 16'd49753, 16'd51831, 16'd15764, 16'd47981, 16'd44120, 16'd61395, 16'd44992, 16'd30740}; // indx = 4478
    #10;
    addra = 32'd143328;
    dina = {96'd0, 16'd49791, 16'd61270, 16'd51784, 16'd56302, 16'd38614, 16'd7509, 16'd17093, 16'd5311, 16'd16466, 16'd11815}; // indx = 4479
    #10;
    addra = 32'd143360;
    dina = {96'd0, 16'd29015, 16'd7126, 16'd62545, 16'd20533, 16'd26012, 16'd47541, 16'd50731, 16'd13750, 16'd2346, 16'd24786}; // indx = 4480
    #10;
    addra = 32'd143392;
    dina = {96'd0, 16'd6691, 16'd18562, 16'd36505, 16'd61375, 16'd39602, 16'd49438, 16'd52237, 16'd59583, 16'd56276, 16'd57420}; // indx = 4481
    #10;
    addra = 32'd143424;
    dina = {96'd0, 16'd14024, 16'd11881, 16'd59257, 16'd26041, 16'd58327, 16'd58562, 16'd62260, 16'd20532, 16'd7665, 16'd50476}; // indx = 4482
    #10;
    addra = 32'd143456;
    dina = {96'd0, 16'd14961, 16'd23204, 16'd31931, 16'd17861, 16'd40978, 16'd58624, 16'd7842, 16'd31528, 16'd37176, 16'd34804}; // indx = 4483
    #10;
    addra = 32'd143488;
    dina = {96'd0, 16'd17836, 16'd17903, 16'd35419, 16'd45656, 16'd15424, 16'd28288, 16'd55473, 16'd21920, 16'd11377, 16'd6985}; // indx = 4484
    #10;
    addra = 32'd143520;
    dina = {96'd0, 16'd183, 16'd54312, 16'd30059, 16'd695, 16'd34990, 16'd24737, 16'd52907, 16'd63639, 16'd51665, 16'd19401}; // indx = 4485
    #10;
    addra = 32'd143552;
    dina = {96'd0, 16'd33909, 16'd23634, 16'd46790, 16'd63093, 16'd54708, 16'd55521, 16'd5432, 16'd18866, 16'd1525, 16'd12396}; // indx = 4486
    #10;
    addra = 32'd143584;
    dina = {96'd0, 16'd65496, 16'd11326, 16'd57955, 16'd63924, 16'd39021, 16'd39595, 16'd5634, 16'd19681, 16'd42850, 16'd45479}; // indx = 4487
    #10;
    addra = 32'd143616;
    dina = {96'd0, 16'd30688, 16'd57385, 16'd1662, 16'd19441, 16'd52689, 16'd45389, 16'd47962, 16'd65106, 16'd49243, 16'd33646}; // indx = 4488
    #10;
    addra = 32'd143648;
    dina = {96'd0, 16'd19441, 16'd62802, 16'd27153, 16'd65395, 16'd33893, 16'd55892, 16'd38288, 16'd8412, 16'd54743, 16'd16412}; // indx = 4489
    #10;
    addra = 32'd143680;
    dina = {96'd0, 16'd5558, 16'd1989, 16'd16917, 16'd6277, 16'd14573, 16'd20447, 16'd31062, 16'd17516, 16'd24198, 16'd3187}; // indx = 4490
    #10;
    addra = 32'd143712;
    dina = {96'd0, 16'd6170, 16'd44182, 16'd26796, 16'd12379, 16'd9060, 16'd57231, 16'd10807, 16'd43728, 16'd59084, 16'd46612}; // indx = 4491
    #10;
    addra = 32'd143744;
    dina = {96'd0, 16'd63453, 16'd65196, 16'd4984, 16'd61859, 16'd62098, 16'd17538, 16'd34071, 16'd36968, 16'd52647, 16'd54471}; // indx = 4492
    #10;
    addra = 32'd143776;
    dina = {96'd0, 16'd17721, 16'd40617, 16'd55827, 16'd37756, 16'd52993, 16'd55431, 16'd60107, 16'd62352, 16'd6356, 16'd53024}; // indx = 4493
    #10;
    addra = 32'd143808;
    dina = {96'd0, 16'd38638, 16'd53904, 16'd34855, 16'd7725, 16'd4479, 16'd47363, 16'd28781, 16'd5086, 16'd62948, 16'd32954}; // indx = 4494
    #10;
    addra = 32'd143840;
    dina = {96'd0, 16'd41646, 16'd27846, 16'd5240, 16'd12414, 16'd62980, 16'd2332, 16'd42382, 16'd1020, 16'd42854, 16'd23661}; // indx = 4495
    #10;
    addra = 32'd143872;
    dina = {96'd0, 16'd22430, 16'd55245, 16'd36611, 16'd51954, 16'd57823, 16'd63708, 16'd47232, 16'd38059, 16'd22333, 16'd2709}; // indx = 4496
    #10;
    addra = 32'd143904;
    dina = {96'd0, 16'd33540, 16'd22554, 16'd14152, 16'd44929, 16'd26081, 16'd25719, 16'd33700, 16'd13882, 16'd1571, 16'd18007}; // indx = 4497
    #10;
    addra = 32'd143936;
    dina = {96'd0, 16'd24044, 16'd28260, 16'd16752, 16'd50075, 16'd3596, 16'd45257, 16'd42919, 16'd50201, 16'd62501, 16'd10402}; // indx = 4498
    #10;
    addra = 32'd143968;
    dina = {96'd0, 16'd4267, 16'd29030, 16'd26540, 16'd12565, 16'd52244, 16'd16008, 16'd4203, 16'd3965, 16'd51962, 16'd33455}; // indx = 4499
    #10;
    addra = 32'd144000;
    dina = {96'd0, 16'd17753, 16'd8402, 16'd10891, 16'd42016, 16'd26057, 16'd2711, 16'd4871, 16'd46045, 16'd24709, 16'd875}; // indx = 4500
    #10;
    addra = 32'd144032;
    dina = {96'd0, 16'd20750, 16'd47153, 16'd13738, 16'd14021, 16'd55666, 16'd29685, 16'd41411, 16'd4820, 16'd9401, 16'd20781}; // indx = 4501
    #10;
    addra = 32'd144064;
    dina = {96'd0, 16'd17421, 16'd41752, 16'd60734, 16'd43168, 16'd41541, 16'd50575, 16'd30013, 16'd51396, 16'd53448, 16'd6613}; // indx = 4502
    #10;
    addra = 32'd144096;
    dina = {96'd0, 16'd17036, 16'd5600, 16'd36799, 16'd38215, 16'd11980, 16'd27506, 16'd37475, 16'd51023, 16'd5655, 16'd33258}; // indx = 4503
    #10;
    addra = 32'd144128;
    dina = {96'd0, 16'd46246, 16'd49051, 16'd3415, 16'd2625, 16'd26346, 16'd64448, 16'd56708, 16'd51685, 16'd18493, 16'd44650}; // indx = 4504
    #10;
    addra = 32'd144160;
    dina = {96'd0, 16'd62336, 16'd24772, 16'd12103, 16'd34314, 16'd6469, 16'd42943, 16'd7115, 16'd7380, 16'd56896, 16'd50551}; // indx = 4505
    #10;
    addra = 32'd144192;
    dina = {96'd0, 16'd44474, 16'd45170, 16'd62473, 16'd54049, 16'd54257, 16'd23086, 16'd32530, 16'd49761, 16'd21959, 16'd20434}; // indx = 4506
    #10;
    addra = 32'd144224;
    dina = {96'd0, 16'd58345, 16'd38249, 16'd16751, 16'd14593, 16'd11261, 16'd48443, 16'd17810, 16'd41405, 16'd6384, 16'd19396}; // indx = 4507
    #10;
    addra = 32'd144256;
    dina = {96'd0, 16'd26714, 16'd34621, 16'd1445, 16'd41519, 16'd45166, 16'd8905, 16'd32906, 16'd11754, 16'd37274, 16'd36679}; // indx = 4508
    #10;
    addra = 32'd144288;
    dina = {96'd0, 16'd10955, 16'd36654, 16'd52944, 16'd48475, 16'd31680, 16'd50620, 16'd3053, 16'd7878, 16'd59178, 16'd6181}; // indx = 4509
    #10;
    addra = 32'd144320;
    dina = {96'd0, 16'd1136, 16'd55215, 16'd40340, 16'd51489, 16'd27133, 16'd20963, 16'd4031, 16'd25805, 16'd49858, 16'd62570}; // indx = 4510
    #10;
    addra = 32'd144352;
    dina = {96'd0, 16'd59569, 16'd9604, 16'd9360, 16'd27796, 16'd465, 16'd9515, 16'd19594, 16'd23651, 16'd6394, 16'd33122}; // indx = 4511
    #10;
    addra = 32'd144384;
    dina = {96'd0, 16'd12827, 16'd54077, 16'd32969, 16'd48853, 16'd11964, 16'd44895, 16'd26195, 16'd56981, 16'd42716, 16'd40614}; // indx = 4512
    #10;
    addra = 32'd144416;
    dina = {96'd0, 16'd57438, 16'd10151, 16'd28910, 16'd22930, 16'd59802, 16'd27606, 16'd26561, 16'd45874, 16'd32974, 16'd22388}; // indx = 4513
    #10;
    addra = 32'd144448;
    dina = {96'd0, 16'd4313, 16'd1535, 16'd45193, 16'd22044, 16'd54008, 16'd12121, 16'd10831, 16'd11084, 16'd36681, 16'd26560}; // indx = 4514
    #10;
    addra = 32'd144480;
    dina = {96'd0, 16'd43813, 16'd202, 16'd10526, 16'd51546, 16'd16841, 16'd5473, 16'd57465, 16'd14121, 16'd35148, 16'd51933}; // indx = 4515
    #10;
    addra = 32'd144512;
    dina = {96'd0, 16'd10197, 16'd41829, 16'd4856, 16'd26252, 16'd36379, 16'd39337, 16'd64937, 16'd43739, 16'd14242, 16'd58651}; // indx = 4516
    #10;
    addra = 32'd144544;
    dina = {96'd0, 16'd38983, 16'd36307, 16'd33210, 16'd5386, 16'd56630, 16'd18228, 16'd30951, 16'd58524, 16'd54615, 16'd26556}; // indx = 4517
    #10;
    addra = 32'd144576;
    dina = {96'd0, 16'd34754, 16'd22414, 16'd20834, 16'd3975, 16'd44866, 16'd10518, 16'd58684, 16'd43468, 16'd48916, 16'd17145}; // indx = 4518
    #10;
    addra = 32'd144608;
    dina = {96'd0, 16'd1982, 16'd8073, 16'd43504, 16'd48582, 16'd8683, 16'd64846, 16'd65297, 16'd27483, 16'd57716, 16'd47409}; // indx = 4519
    #10;
    addra = 32'd144640;
    dina = {96'd0, 16'd51547, 16'd41325, 16'd46408, 16'd15236, 16'd63279, 16'd8243, 16'd11760, 16'd1180, 16'd5667, 16'd35808}; // indx = 4520
    #10;
    addra = 32'd144672;
    dina = {96'd0, 16'd65181, 16'd36830, 16'd63368, 16'd16120, 16'd28494, 16'd1478, 16'd9925, 16'd10452, 16'd57466, 16'd9313}; // indx = 4521
    #10;
    addra = 32'd144704;
    dina = {96'd0, 16'd55429, 16'd45401, 16'd10223, 16'd39969, 16'd63967, 16'd29194, 16'd38756, 16'd18513, 16'd7412, 16'd63759}; // indx = 4522
    #10;
    addra = 32'd144736;
    dina = {96'd0, 16'd26225, 16'd64351, 16'd16251, 16'd63350, 16'd58004, 16'd22771, 16'd8239, 16'd1806, 16'd61580, 16'd52249}; // indx = 4523
    #10;
    addra = 32'd144768;
    dina = {96'd0, 16'd48793, 16'd62544, 16'd30374, 16'd47903, 16'd22535, 16'd55692, 16'd41786, 16'd16950, 16'd25280, 16'd2162}; // indx = 4524
    #10;
    addra = 32'd144800;
    dina = {96'd0, 16'd32998, 16'd59043, 16'd18021, 16'd33477, 16'd53296, 16'd24586, 16'd7149, 16'd13096, 16'd60584, 16'd9997}; // indx = 4525
    #10;
    addra = 32'd144832;
    dina = {96'd0, 16'd17150, 16'd7389, 16'd61585, 16'd62602, 16'd42294, 16'd52198, 16'd63326, 16'd50766, 16'd2368, 16'd59844}; // indx = 4526
    #10;
    addra = 32'd144864;
    dina = {96'd0, 16'd53064, 16'd54554, 16'd47334, 16'd8671, 16'd24328, 16'd46480, 16'd33061, 16'd14448, 16'd20711, 16'd63595}; // indx = 4527
    #10;
    addra = 32'd144896;
    dina = {96'd0, 16'd49171, 16'd34908, 16'd16788, 16'd62673, 16'd16805, 16'd27644, 16'd45990, 16'd25568, 16'd64842, 16'd40912}; // indx = 4528
    #10;
    addra = 32'd144928;
    dina = {96'd0, 16'd20573, 16'd61061, 16'd48343, 16'd19194, 16'd60784, 16'd45165, 16'd20196, 16'd62287, 16'd45673, 16'd29856}; // indx = 4529
    #10;
    addra = 32'd144960;
    dina = {96'd0, 16'd32115, 16'd49016, 16'd57546, 16'd49005, 16'd24091, 16'd48526, 16'd11430, 16'd25790, 16'd61996, 16'd6905}; // indx = 4530
    #10;
    addra = 32'd144992;
    dina = {96'd0, 16'd7748, 16'd6539, 16'd48939, 16'd12470, 16'd35291, 16'd3034, 16'd44609, 16'd5436, 16'd32052, 16'd23664}; // indx = 4531
    #10;
    addra = 32'd145024;
    dina = {96'd0, 16'd6014, 16'd53558, 16'd21064, 16'd44999, 16'd52994, 16'd17248, 16'd30973, 16'd37974, 16'd682, 16'd22735}; // indx = 4532
    #10;
    addra = 32'd145056;
    dina = {96'd0, 16'd49894, 16'd36673, 16'd60664, 16'd25238, 16'd39239, 16'd33001, 16'd27675, 16'd53622, 16'd14953, 16'd53162}; // indx = 4533
    #10;
    addra = 32'd145088;
    dina = {96'd0, 16'd28158, 16'd10274, 16'd39560, 16'd17713, 16'd43767, 16'd13082, 16'd63289, 16'd27669, 16'd26961, 16'd57464}; // indx = 4534
    #10;
    addra = 32'd145120;
    dina = {96'd0, 16'd60658, 16'd39727, 16'd31700, 16'd12409, 16'd41364, 16'd17332, 16'd29839, 16'd48020, 16'd13671, 16'd47369}; // indx = 4535
    #10;
    addra = 32'd145152;
    dina = {96'd0, 16'd8020, 16'd45928, 16'd60085, 16'd48331, 16'd52646, 16'd38580, 16'd23339, 16'd40229, 16'd56066, 16'd21557}; // indx = 4536
    #10;
    addra = 32'd145184;
    dina = {96'd0, 16'd26742, 16'd10947, 16'd64057, 16'd21045, 16'd3208, 16'd239, 16'd59147, 16'd9341, 16'd45740, 16'd24730}; // indx = 4537
    #10;
    addra = 32'd145216;
    dina = {96'd0, 16'd20247, 16'd56719, 16'd54712, 16'd7959, 16'd17789, 16'd21009, 16'd52106, 16'd43955, 16'd59144, 16'd36685}; // indx = 4538
    #10;
    addra = 32'd145248;
    dina = {96'd0, 16'd4900, 16'd59812, 16'd63776, 16'd2947, 16'd7015, 16'd44955, 16'd18080, 16'd50279, 16'd51317, 16'd16232}; // indx = 4539
    #10;
    addra = 32'd145280;
    dina = {96'd0, 16'd31067, 16'd24699, 16'd57874, 16'd47920, 16'd29886, 16'd3579, 16'd51838, 16'd6536, 16'd35583, 16'd46697}; // indx = 4540
    #10;
    addra = 32'd145312;
    dina = {96'd0, 16'd11473, 16'd23771, 16'd24121, 16'd49641, 16'd19829, 16'd29225, 16'd61188, 16'd33884, 16'd45586, 16'd26366}; // indx = 4541
    #10;
    addra = 32'd145344;
    dina = {96'd0, 16'd60545, 16'd48567, 16'd326, 16'd61680, 16'd39889, 16'd57862, 16'd46514, 16'd64496, 16'd270, 16'd45124}; // indx = 4542
    #10;
    addra = 32'd145376;
    dina = {96'd0, 16'd53260, 16'd34259, 16'd47616, 16'd45659, 16'd62218, 16'd60175, 16'd27511, 16'd44050, 16'd15007, 16'd38672}; // indx = 4543
    #10;
    addra = 32'd145408;
    dina = {96'd0, 16'd27833, 16'd4017, 16'd909, 16'd41330, 16'd54245, 16'd29237, 16'd32532, 16'd274, 16'd3938, 16'd7905}; // indx = 4544
    #10;
    addra = 32'd145440;
    dina = {96'd0, 16'd14165, 16'd45604, 16'd15231, 16'd12822, 16'd32819, 16'd62852, 16'd13664, 16'd4726, 16'd63342, 16'd42816}; // indx = 4545
    #10;
    addra = 32'd145472;
    dina = {96'd0, 16'd63192, 16'd42198, 16'd34494, 16'd10310, 16'd32885, 16'd22688, 16'd65433, 16'd22595, 16'd36557, 16'd55228}; // indx = 4546
    #10;
    addra = 32'd145504;
    dina = {96'd0, 16'd2069, 16'd40010, 16'd63982, 16'd11490, 16'd41385, 16'd29715, 16'd43114, 16'd44854, 16'd10972, 16'd53789}; // indx = 4547
    #10;
    addra = 32'd145536;
    dina = {96'd0, 16'd61601, 16'd25936, 16'd73, 16'd23104, 16'd48270, 16'd23284, 16'd3924, 16'd38707, 16'd21974, 16'd4277}; // indx = 4548
    #10;
    addra = 32'd145568;
    dina = {96'd0, 16'd22655, 16'd34359, 16'd14790, 16'd41254, 16'd55763, 16'd11648, 16'd51105, 16'd40878, 16'd14142, 16'd27540}; // indx = 4549
    #10;
    addra = 32'd145600;
    dina = {96'd0, 16'd20711, 16'd63826, 16'd62419, 16'd5280, 16'd44215, 16'd53064, 16'd623, 16'd7332, 16'd692, 16'd1119}; // indx = 4550
    #10;
    addra = 32'd145632;
    dina = {96'd0, 16'd58953, 16'd57674, 16'd57067, 16'd43620, 16'd43299, 16'd52690, 16'd39201, 16'd37144, 16'd65090, 16'd3749}; // indx = 4551
    #10;
    addra = 32'd145664;
    dina = {96'd0, 16'd32806, 16'd29700, 16'd22178, 16'd34236, 16'd49531, 16'd57280, 16'd24108, 16'd16632, 16'd11413, 16'd47052}; // indx = 4552
    #10;
    addra = 32'd145696;
    dina = {96'd0, 16'd40511, 16'd30583, 16'd45588, 16'd35641, 16'd18010, 16'd46983, 16'd42365, 16'd50248, 16'd5764, 16'd4210}; // indx = 4553
    #10;
    addra = 32'd145728;
    dina = {96'd0, 16'd45179, 16'd40626, 16'd62762, 16'd52054, 16'd47561, 16'd41501, 16'd14404, 16'd21240, 16'd55075, 16'd60603}; // indx = 4554
    #10;
    addra = 32'd145760;
    dina = {96'd0, 16'd48163, 16'd26116, 16'd5963, 16'd53970, 16'd34879, 16'd33666, 16'd39438, 16'd26523, 16'd28533, 16'd62372}; // indx = 4555
    #10;
    addra = 32'd145792;
    dina = {96'd0, 16'd7065, 16'd59587, 16'd62699, 16'd10990, 16'd55228, 16'd9837, 16'd23700, 16'd5858, 16'd26507, 16'd334}; // indx = 4556
    #10;
    addra = 32'd145824;
    dina = {96'd0, 16'd34002, 16'd46228, 16'd37047, 16'd32359, 16'd50918, 16'd63300, 16'd31045, 16'd39087, 16'd46858, 16'd21460}; // indx = 4557
    #10;
    addra = 32'd145856;
    dina = {96'd0, 16'd1668, 16'd42030, 16'd46443, 16'd38217, 16'd60868, 16'd49348, 16'd28201, 16'd22488, 16'd53219, 16'd8095}; // indx = 4558
    #10;
    addra = 32'd145888;
    dina = {96'd0, 16'd9644, 16'd14946, 16'd50514, 16'd28757, 16'd21384, 16'd36882, 16'd61505, 16'd62564, 16'd21451, 16'd25659}; // indx = 4559
    #10;
    addra = 32'd145920;
    dina = {96'd0, 16'd31321, 16'd12859, 16'd4795, 16'd26953, 16'd26817, 16'd22907, 16'd1748, 16'd49416, 16'd1023, 16'd2207}; // indx = 4560
    #10;
    addra = 32'd145952;
    dina = {96'd0, 16'd52131, 16'd65223, 16'd34660, 16'd28610, 16'd34973, 16'd31756, 16'd11761, 16'd58742, 16'd41194, 16'd57329}; // indx = 4561
    #10;
    addra = 32'd145984;
    dina = {96'd0, 16'd14103, 16'd53610, 16'd46727, 16'd60977, 16'd10314, 16'd29759, 16'd60838, 16'd7879, 16'd5223, 16'd19501}; // indx = 4562
    #10;
    addra = 32'd146016;
    dina = {96'd0, 16'd54483, 16'd32690, 16'd46736, 16'd34194, 16'd11383, 16'd57726, 16'd21881, 16'd49948, 16'd23649, 16'd41209}; // indx = 4563
    #10;
    addra = 32'd146048;
    dina = {96'd0, 16'd48149, 16'd10557, 16'd53011, 16'd17427, 16'd44809, 16'd50462, 16'd47546, 16'd24722, 16'd24072, 16'd49663}; // indx = 4564
    #10;
    addra = 32'd146080;
    dina = {96'd0, 16'd6989, 16'd13735, 16'd29814, 16'd23329, 16'd57938, 16'd51662, 16'd37064, 16'd24219, 16'd44206, 16'd44696}; // indx = 4565
    #10;
    addra = 32'd146112;
    dina = {96'd0, 16'd57292, 16'd11436, 16'd1840, 16'd30122, 16'd15406, 16'd2175, 16'd39420, 16'd28443, 16'd23656, 16'd19418}; // indx = 4566
    #10;
    addra = 32'd146144;
    dina = {96'd0, 16'd11475, 16'd24050, 16'd50686, 16'd48608, 16'd11127, 16'd46912, 16'd19818, 16'd12117, 16'd46121, 16'd57830}; // indx = 4567
    #10;
    addra = 32'd146176;
    dina = {96'd0, 16'd13681, 16'd19766, 16'd47297, 16'd38347, 16'd57259, 16'd13762, 16'd27742, 16'd16540, 16'd10571, 16'd51154}; // indx = 4568
    #10;
    addra = 32'd146208;
    dina = {96'd0, 16'd40445, 16'd12781, 16'd33104, 16'd26017, 16'd7381, 16'd23586, 16'd46053, 16'd32324, 16'd50802, 16'd8145}; // indx = 4569
    #10;
    addra = 32'd146240;
    dina = {96'd0, 16'd63740, 16'd57593, 16'd43939, 16'd18859, 16'd33970, 16'd44496, 16'd49157, 16'd292, 16'd53177, 16'd57667}; // indx = 4570
    #10;
    addra = 32'd146272;
    dina = {96'd0, 16'd28711, 16'd58425, 16'd47224, 16'd42694, 16'd17302, 16'd45510, 16'd27436, 16'd27746, 16'd28387, 16'd23877}; // indx = 4571
    #10;
    addra = 32'd146304;
    dina = {96'd0, 16'd54565, 16'd23828, 16'd41996, 16'd57427, 16'd19697, 16'd62507, 16'd42679, 16'd52596, 16'd45304, 16'd65104}; // indx = 4572
    #10;
    addra = 32'd146336;
    dina = {96'd0, 16'd13821, 16'd33542, 16'd47636, 16'd64111, 16'd43695, 16'd38347, 16'd32041, 16'd40043, 16'd5139, 16'd36349}; // indx = 4573
    #10;
    addra = 32'd146368;
    dina = {96'd0, 16'd61448, 16'd46111, 16'd20347, 16'd15693, 16'd51465, 16'd35131, 16'd46270, 16'd21630, 16'd43672, 16'd30731}; // indx = 4574
    #10;
    addra = 32'd146400;
    dina = {96'd0, 16'd21071, 16'd164, 16'd25570, 16'd49583, 16'd10195, 16'd35441, 16'd49442, 16'd53071, 16'd3293, 16'd2444}; // indx = 4575
    #10;
    addra = 32'd146432;
    dina = {96'd0, 16'd4714, 16'd39098, 16'd19261, 16'd40096, 16'd5053, 16'd36063, 16'd9188, 16'd57404, 16'd37371, 16'd48300}; // indx = 4576
    #10;
    addra = 32'd146464;
    dina = {96'd0, 16'd4424, 16'd25883, 16'd21644, 16'd2218, 16'd59375, 16'd18325, 16'd27662, 16'd25758, 16'd46764, 16'd59805}; // indx = 4577
    #10;
    addra = 32'd146496;
    dina = {96'd0, 16'd60610, 16'd36255, 16'd65105, 16'd46999, 16'd44653, 16'd60979, 16'd4678, 16'd55172, 16'd40620, 16'd23927}; // indx = 4578
    #10;
    addra = 32'd146528;
    dina = {96'd0, 16'd47391, 16'd45725, 16'd50285, 16'd33811, 16'd30742, 16'd14096, 16'd37191, 16'd48784, 16'd14625, 16'd589}; // indx = 4579
    #10;
    addra = 32'd146560;
    dina = {96'd0, 16'd62577, 16'd41489, 16'd24191, 16'd28920, 16'd50229, 16'd16574, 16'd65476, 16'd6071, 16'd17112, 16'd50621}; // indx = 4580
    #10;
    addra = 32'd146592;
    dina = {96'd0, 16'd30861, 16'd32405, 16'd18854, 16'd54755, 16'd16419, 16'd27637, 16'd51597, 16'd3054, 16'd53336, 16'd9246}; // indx = 4581
    #10;
    addra = 32'd146624;
    dina = {96'd0, 16'd5533, 16'd38116, 16'd23788, 16'd49071, 16'd31723, 16'd20082, 16'd64113, 16'd1743, 16'd56874, 16'd40837}; // indx = 4582
    #10;
    addra = 32'd146656;
    dina = {96'd0, 16'd44482, 16'd16144, 16'd58602, 16'd338, 16'd45380, 16'd9937, 16'd358, 16'd52846, 16'd10607, 16'd45746}; // indx = 4583
    #10;
    addra = 32'd146688;
    dina = {96'd0, 16'd76, 16'd21039, 16'd45970, 16'd3797, 16'd17367, 16'd50902, 16'd27045, 16'd34269, 16'd34402, 16'd41523}; // indx = 4584
    #10;
    addra = 32'd146720;
    dina = {96'd0, 16'd59897, 16'd48351, 16'd3238, 16'd31462, 16'd38080, 16'd56235, 16'd59329, 16'd59296, 16'd44802, 16'd9416}; // indx = 4585
    #10;
    addra = 32'd146752;
    dina = {96'd0, 16'd47763, 16'd60636, 16'd2444, 16'd16697, 16'd46696, 16'd53114, 16'd29861, 16'd23713, 16'd51675, 16'd64111}; // indx = 4586
    #10;
    addra = 32'd146784;
    dina = {96'd0, 16'd25040, 16'd28927, 16'd6637, 16'd63541, 16'd1197, 16'd52328, 16'd4336, 16'd37041, 16'd45928, 16'd13058}; // indx = 4587
    #10;
    addra = 32'd146816;
    dina = {96'd0, 16'd4351, 16'd60050, 16'd43325, 16'd26232, 16'd60504, 16'd58035, 16'd25486, 16'd35446, 16'd42215, 16'd1480}; // indx = 4588
    #10;
    addra = 32'd146848;
    dina = {96'd0, 16'd43368, 16'd5510, 16'd54648, 16'd9240, 16'd59182, 16'd37102, 16'd24212, 16'd36840, 16'd8747, 16'd49267}; // indx = 4589
    #10;
    addra = 32'd146880;
    dina = {96'd0, 16'd40013, 16'd21042, 16'd14011, 16'd4120, 16'd60033, 16'd35080, 16'd34250, 16'd40047, 16'd59554, 16'd6830}; // indx = 4590
    #10;
    addra = 32'd146912;
    dina = {96'd0, 16'd57992, 16'd49843, 16'd43299, 16'd21576, 16'd39554, 16'd20616, 16'd18141, 16'd30814, 16'd14837, 16'd8833}; // indx = 4591
    #10;
    addra = 32'd146944;
    dina = {96'd0, 16'd54758, 16'd44925, 16'd31067, 16'd46746, 16'd35013, 16'd20236, 16'd55435, 16'd64538, 16'd47596, 16'd12332}; // indx = 4592
    #10;
    addra = 32'd146976;
    dina = {96'd0, 16'd19160, 16'd36562, 16'd37769, 16'd47876, 16'd699, 16'd43636, 16'd1514, 16'd31561, 16'd49048, 16'd44298}; // indx = 4593
    #10;
    addra = 32'd147008;
    dina = {96'd0, 16'd45885, 16'd24017, 16'd30801, 16'd62336, 16'd8883, 16'd920, 16'd34443, 16'd28049, 16'd16517, 16'd61728}; // indx = 4594
    #10;
    addra = 32'd147040;
    dina = {96'd0, 16'd29655, 16'd12905, 16'd61929, 16'd14136, 16'd54850, 16'd44607, 16'd51225, 16'd37859, 16'd39675, 16'd3899}; // indx = 4595
    #10;
    addra = 32'd147072;
    dina = {96'd0, 16'd64383, 16'd9124, 16'd52227, 16'd4001, 16'd55371, 16'd2778, 16'd29087, 16'd35822, 16'd33086, 16'd36268}; // indx = 4596
    #10;
    addra = 32'd147104;
    dina = {96'd0, 16'd19481, 16'd45288, 16'd43398, 16'd46782, 16'd60960, 16'd49908, 16'd24759, 16'd21639, 16'd37874, 16'd59820}; // indx = 4597
    #10;
    addra = 32'd147136;
    dina = {96'd0, 16'd16811, 16'd55521, 16'd38788, 16'd30866, 16'd40279, 16'd37088, 16'd51000, 16'd10067, 16'd7750, 16'd7893}; // indx = 4598
    #10;
    addra = 32'd147168;
    dina = {96'd0, 16'd28399, 16'd19686, 16'd30449, 16'd28132, 16'd16639, 16'd18641, 16'd55431, 16'd58942, 16'd60609, 16'd61496}; // indx = 4599
    #10;
    addra = 32'd147200;
    dina = {96'd0, 16'd34283, 16'd7975, 16'd39827, 16'd53426, 16'd40769, 16'd8577, 16'd36105, 16'd43975, 16'd28534, 16'd13154}; // indx = 4600
    #10;
    addra = 32'd147232;
    dina = {96'd0, 16'd35494, 16'd29361, 16'd23153, 16'd22490, 16'd10114, 16'd49564, 16'd55240, 16'd35398, 16'd43715, 16'd56358}; // indx = 4601
    #10;
    addra = 32'd147264;
    dina = {96'd0, 16'd26374, 16'd63257, 16'd23049, 16'd26134, 16'd16987, 16'd46732, 16'd10210, 16'd62586, 16'd43147, 16'd62107}; // indx = 4602
    #10;
    addra = 32'd147296;
    dina = {96'd0, 16'd2080, 16'd26755, 16'd47759, 16'd61836, 16'd16234, 16'd60769, 16'd996, 16'd17495, 16'd27397, 16'd32873}; // indx = 4603
    #10;
    addra = 32'd147328;
    dina = {96'd0, 16'd22154, 16'd56739, 16'd11596, 16'd54158, 16'd13445, 16'd52788, 16'd27244, 16'd39724, 16'd64805, 16'd20811}; // indx = 4604
    #10;
    addra = 32'd147360;
    dina = {96'd0, 16'd63546, 16'd53013, 16'd64408, 16'd24930, 16'd21632, 16'd43803, 16'd3176, 16'd40047, 16'd148, 16'd12264}; // indx = 4605
    #10;
    addra = 32'd147392;
    dina = {96'd0, 16'd18678, 16'd59673, 16'd62671, 16'd11417, 16'd40909, 16'd24689, 16'd23002, 16'd16818, 16'd32481, 16'd14968}; // indx = 4606
    #10;
    addra = 32'd147424;
    dina = {96'd0, 16'd44483, 16'd50715, 16'd49410, 16'd60027, 16'd38545, 16'd16085, 16'd18567, 16'd46233, 16'd10461, 16'd44946}; // indx = 4607
    #10;
    addra = 32'd147456;
    dina = {96'd0, 16'd4461, 16'd25247, 16'd40400, 16'd48251, 16'd34463, 16'd11915, 16'd5713, 16'd13917, 16'd27151, 16'd16390}; // indx = 4608
    #10;
    addra = 32'd147488;
    dina = {96'd0, 16'd59606, 16'd34822, 16'd30538, 16'd40605, 16'd42336, 16'd44457, 16'd42920, 16'd60213, 16'd16445, 16'd1858}; // indx = 4609
    #10;
    addra = 32'd147520;
    dina = {96'd0, 16'd8294, 16'd42853, 16'd16585, 16'd39184, 16'd40406, 16'd20381, 16'd35902, 16'd12784, 16'd45396, 16'd49897}; // indx = 4610
    #10;
    addra = 32'd147552;
    dina = {96'd0, 16'd24795, 16'd35758, 16'd59748, 16'd22849, 16'd4934, 16'd49882, 16'd19563, 16'd17363, 16'd11217, 16'd3160}; // indx = 4611
    #10;
    addra = 32'd147584;
    dina = {96'd0, 16'd61506, 16'd5120, 16'd44217, 16'd46071, 16'd31261, 16'd21856, 16'd24927, 16'd35194, 16'd64431, 16'd35896}; // indx = 4612
    #10;
    addra = 32'd147616;
    dina = {96'd0, 16'd40634, 16'd65302, 16'd971, 16'd5490, 16'd38439, 16'd17846, 16'd2165, 16'd64618, 16'd20587, 16'd28488}; // indx = 4613
    #10;
    addra = 32'd147648;
    dina = {96'd0, 16'd57906, 16'd59483, 16'd62132, 16'd33902, 16'd1786, 16'd56655, 16'd11707, 16'd13523, 16'd14225, 16'd33608}; // indx = 4614
    #10;
    addra = 32'd147680;
    dina = {96'd0, 16'd40270, 16'd9104, 16'd50077, 16'd12096, 16'd8798, 16'd30015, 16'd11723, 16'd48936, 16'd61940, 16'd54690}; // indx = 4615
    #10;
    addra = 32'd147712;
    dina = {96'd0, 16'd40239, 16'd17816, 16'd35382, 16'd47300, 16'd38802, 16'd7973, 16'd51226, 16'd18631, 16'd24841, 16'd40899}; // indx = 4616
    #10;
    addra = 32'd147744;
    dina = {96'd0, 16'd19262, 16'd28000, 16'd24314, 16'd14727, 16'd57182, 16'd6566, 16'd36310, 16'd28124, 16'd63837, 16'd61512}; // indx = 4617
    #10;
    addra = 32'd147776;
    dina = {96'd0, 16'd28076, 16'd61135, 16'd9412, 16'd2231, 16'd26675, 16'd39317, 16'd2459, 16'd24406, 16'd10867, 16'd59471}; // indx = 4618
    #10;
    addra = 32'd147808;
    dina = {96'd0, 16'd35162, 16'd27749, 16'd30888, 16'd38028, 16'd4600, 16'd50326, 16'd16944, 16'd10997, 16'd44847, 16'd54619}; // indx = 4619
    #10;
    addra = 32'd147840;
    dina = {96'd0, 16'd29457, 16'd10273, 16'd51138, 16'd10039, 16'd9943, 16'd37993, 16'd63449, 16'd8802, 16'd54948, 16'd6711}; // indx = 4620
    #10;
    addra = 32'd147872;
    dina = {96'd0, 16'd32009, 16'd21370, 16'd47291, 16'd6794, 16'd62926, 16'd22282, 16'd45370, 16'd43015, 16'd24550, 16'd30718}; // indx = 4621
    #10;
    addra = 32'd147904;
    dina = {96'd0, 16'd28778, 16'd57652, 16'd11782, 16'd24966, 16'd18102, 16'd12609, 16'd48069, 16'd33392, 16'd23374, 16'd6472}; // indx = 4622
    #10;
    addra = 32'd147936;
    dina = {96'd0, 16'd13800, 16'd46414, 16'd21124, 16'd2391, 16'd44860, 16'd64052, 16'd50026, 16'd31131, 16'd39418, 16'd27192}; // indx = 4623
    #10;
    addra = 32'd147968;
    dina = {96'd0, 16'd11445, 16'd2970, 16'd46563, 16'd48670, 16'd34572, 16'd3919, 16'd21710, 16'd9141, 16'd368, 16'd36063}; // indx = 4624
    #10;
    addra = 32'd148000;
    dina = {96'd0, 16'd46896, 16'd11207, 16'd5522, 16'd49846, 16'd16664, 16'd17887, 16'd30342, 16'd64139, 16'd46602, 16'd8462}; // indx = 4625
    #10;
    addra = 32'd148032;
    dina = {96'd0, 16'd48284, 16'd57721, 16'd51881, 16'd21040, 16'd24490, 16'd8966, 16'd12742, 16'd20491, 16'd53171, 16'd602}; // indx = 4626
    #10;
    addra = 32'd148064;
    dina = {96'd0, 16'd14486, 16'd12625, 16'd52232, 16'd16359, 16'd21283, 16'd17875, 16'd36895, 16'd1638, 16'd1168, 16'd4374}; // indx = 4627
    #10;
    addra = 32'd148096;
    dina = {96'd0, 16'd38027, 16'd41046, 16'd45776, 16'd22889, 16'd15672, 16'd19860, 16'd23921, 16'd762, 16'd21938, 16'd29874}; // indx = 4628
    #10;
    addra = 32'd148128;
    dina = {96'd0, 16'd12599, 16'd53761, 16'd3170, 16'd63244, 16'd55222, 16'd8471, 16'd44255, 16'd32208, 16'd43657, 16'd39511}; // indx = 4629
    #10;
    addra = 32'd148160;
    dina = {96'd0, 16'd31613, 16'd62312, 16'd64311, 16'd59619, 16'd6729, 16'd63242, 16'd45654, 16'd23548, 16'd63165, 16'd39068}; // indx = 4630
    #10;
    addra = 32'd148192;
    dina = {96'd0, 16'd7163, 16'd17512, 16'd8554, 16'd61182, 16'd14398, 16'd39500, 16'd47182, 16'd29669, 16'd27258, 16'd28978}; // indx = 4631
    #10;
    addra = 32'd148224;
    dina = {96'd0, 16'd57848, 16'd23807, 16'd1541, 16'd21962, 16'd29110, 16'd51689, 16'd29532, 16'd6731, 16'd53639, 16'd11975}; // indx = 4632
    #10;
    addra = 32'd148256;
    dina = {96'd0, 16'd57087, 16'd596, 16'd44801, 16'd17872, 16'd17870, 16'd17228, 16'd33485, 16'd62372, 16'd39450, 16'd16133}; // indx = 4633
    #10;
    addra = 32'd148288;
    dina = {96'd0, 16'd2969, 16'd27681, 16'd55305, 16'd20305, 16'd32670, 16'd50924, 16'd63125, 16'd45596, 16'd47777, 16'd4006}; // indx = 4634
    #10;
    addra = 32'd148320;
    dina = {96'd0, 16'd35262, 16'd15438, 16'd39377, 16'd39717, 16'd59429, 16'd50043, 16'd59270, 16'd19095, 16'd57708, 16'd55073}; // indx = 4635
    #10;
    addra = 32'd148352;
    dina = {96'd0, 16'd22563, 16'd4332, 16'd31012, 16'd25903, 16'd42620, 16'd30724, 16'd37136, 16'd41354, 16'd63524, 16'd48158}; // indx = 4636
    #10;
    addra = 32'd148384;
    dina = {96'd0, 16'd55272, 16'd39511, 16'd13000, 16'd28239, 16'd23505, 16'd44389, 16'd63318, 16'd41052, 16'd19846, 16'd56653}; // indx = 4637
    #10;
    addra = 32'd148416;
    dina = {96'd0, 16'd35577, 16'd44205, 16'd63155, 16'd11080, 16'd41141, 16'd57350, 16'd10597, 16'd51209, 16'd60235, 16'd30286}; // indx = 4638
    #10;
    addra = 32'd148448;
    dina = {96'd0, 16'd12182, 16'd10998, 16'd22021, 16'd12819, 16'd9223, 16'd21986, 16'd44501, 16'd7517, 16'd27954, 16'd39081}; // indx = 4639
    #10;
    addra = 32'd148480;
    dina = {96'd0, 16'd53955, 16'd13925, 16'd5017, 16'd24460, 16'd254, 16'd29373, 16'd21936, 16'd6040, 16'd36878, 16'd59957}; // indx = 4640
    #10;
    addra = 32'd148512;
    dina = {96'd0, 16'd30812, 16'd29349, 16'd47084, 16'd22768, 16'd23047, 16'd6132, 16'd31886, 16'd61680, 16'd41218, 16'd44429}; // indx = 4641
    #10;
    addra = 32'd148544;
    dina = {96'd0, 16'd18833, 16'd39217, 16'd4562, 16'd42505, 16'd26181, 16'd11004, 16'd62242, 16'd1416, 16'd60186, 16'd28433}; // indx = 4642
    #10;
    addra = 32'd148576;
    dina = {96'd0, 16'd24119, 16'd62571, 16'd47681, 16'd37979, 16'd58397, 16'd46555, 16'd63496, 16'd21822, 16'd43645, 16'd198}; // indx = 4643
    #10;
    addra = 32'd148608;
    dina = {96'd0, 16'd18884, 16'd46458, 16'd38943, 16'd18122, 16'd46323, 16'd22875, 16'd49403, 16'd36793, 16'd15890, 16'd24886}; // indx = 4644
    #10;
    addra = 32'd148640;
    dina = {96'd0, 16'd41730, 16'd4908, 16'd41247, 16'd60412, 16'd50879, 16'd42753, 16'd63390, 16'd31256, 16'd10904, 16'd50067}; // indx = 4645
    #10;
    addra = 32'd148672;
    dina = {96'd0, 16'd24115, 16'd59730, 16'd55459, 16'd36889, 16'd54926, 16'd47808, 16'd52037, 16'd2286, 16'd2229, 16'd59236}; // indx = 4646
    #10;
    addra = 32'd148704;
    dina = {96'd0, 16'd6677, 16'd33824, 16'd61877, 16'd3710, 16'd24951, 16'd5227, 16'd38793, 16'd57732, 16'd36098, 16'd27859}; // indx = 4647
    #10;
    addra = 32'd148736;
    dina = {96'd0, 16'd26892, 16'd45150, 16'd64229, 16'd9186, 16'd41328, 16'd23943, 16'd539, 16'd18655, 16'd2864, 16'd45366}; // indx = 4648
    #10;
    addra = 32'd148768;
    dina = {96'd0, 16'd19160, 16'd25777, 16'd15824, 16'd30162, 16'd22599, 16'd48794, 16'd64709, 16'd4663, 16'd1601, 16'd41363}; // indx = 4649
    #10;
    addra = 32'd148800;
    dina = {96'd0, 16'd6417, 16'd38901, 16'd26777, 16'd38581, 16'd27514, 16'd18221, 16'd22131, 16'd36384, 16'd58450, 16'd15724}; // indx = 4650
    #10;
    addra = 32'd148832;
    dina = {96'd0, 16'd39035, 16'd49640, 16'd35786, 16'd37712, 16'd65389, 16'd15081, 16'd48741, 16'd1026, 16'd16288, 16'd45192}; // indx = 4651
    #10;
    addra = 32'd148864;
    dina = {96'd0, 16'd49040, 16'd53236, 16'd31434, 16'd13659, 16'd30954, 16'd7314, 16'd46098, 16'd24867, 16'd51406, 16'd22680}; // indx = 4652
    #10;
    addra = 32'd148896;
    dina = {96'd0, 16'd61615, 16'd65251, 16'd47834, 16'd45698, 16'd38290, 16'd12160, 16'd42313, 16'd54865, 16'd30266, 16'd3604}; // indx = 4653
    #10;
    addra = 32'd148928;
    dina = {96'd0, 16'd11322, 16'd18450, 16'd48947, 16'd9357, 16'd57452, 16'd15059, 16'd41636, 16'd24782, 16'd43749, 16'd23701}; // indx = 4654
    #10;
    addra = 32'd148960;
    dina = {96'd0, 16'd19086, 16'd35245, 16'd58229, 16'd13757, 16'd18147, 16'd59887, 16'd9114, 16'd25528, 16'd20109, 16'd23245}; // indx = 4655
    #10;
    addra = 32'd148992;
    dina = {96'd0, 16'd28737, 16'd61548, 16'd18898, 16'd24361, 16'd23686, 16'd25528, 16'd58534, 16'd30811, 16'd12910, 16'd21848}; // indx = 4656
    #10;
    addra = 32'd149024;
    dina = {96'd0, 16'd55849, 16'd51204, 16'd56747, 16'd62536, 16'd53498, 16'd16806, 16'd43767, 16'd18628, 16'd58374, 16'd58204}; // indx = 4657
    #10;
    addra = 32'd149056;
    dina = {96'd0, 16'd46240, 16'd13720, 16'd61788, 16'd36176, 16'd13601, 16'd10865, 16'd4104, 16'd913, 16'd11644, 16'd31871}; // indx = 4658
    #10;
    addra = 32'd149088;
    dina = {96'd0, 16'd1321, 16'd41345, 16'd27027, 16'd28605, 16'd54282, 16'd21520, 16'd48311, 16'd40082, 16'd51101, 16'd30999}; // indx = 4659
    #10;
    addra = 32'd149120;
    dina = {96'd0, 16'd14212, 16'd53236, 16'd6236, 16'd50732, 16'd39426, 16'd5321, 16'd20991, 16'd25957, 16'd53678, 16'd8855}; // indx = 4660
    #10;
    addra = 32'd149152;
    dina = {96'd0, 16'd23072, 16'd37674, 16'd30236, 16'd31546, 16'd57956, 16'd65030, 16'd23934, 16'd44299, 16'd2339, 16'd38532}; // indx = 4661
    #10;
    addra = 32'd149184;
    dina = {96'd0, 16'd12374, 16'd22329, 16'd33556, 16'd57446, 16'd17506, 16'd895, 16'd25175, 16'd39644, 16'd48520, 16'd31406}; // indx = 4662
    #10;
    addra = 32'd149216;
    dina = {96'd0, 16'd341, 16'd17892, 16'd59699, 16'd53976, 16'd11589, 16'd48785, 16'd7074, 16'd19706, 16'd9437, 16'd61349}; // indx = 4663
    #10;
    addra = 32'd149248;
    dina = {96'd0, 16'd19558, 16'd63941, 16'd47117, 16'd25291, 16'd53463, 16'd8664, 16'd15532, 16'd31241, 16'd902, 16'd36791}; // indx = 4664
    #10;
    addra = 32'd149280;
    dina = {96'd0, 16'd29854, 16'd53979, 16'd10945, 16'd60008, 16'd966, 16'd22529, 16'd30541, 16'd34747, 16'd33887, 16'd38567}; // indx = 4665
    #10;
    addra = 32'd149312;
    dina = {96'd0, 16'd24373, 16'd46117, 16'd42156, 16'd1432, 16'd19888, 16'd33141, 16'd20112, 16'd11720, 16'd47739, 16'd35887}; // indx = 4666
    #10;
    addra = 32'd149344;
    dina = {96'd0, 16'd22473, 16'd16876, 16'd8830, 16'd7583, 16'd16441, 16'd21185, 16'd9410, 16'd40135, 16'd15963, 16'd51005}; // indx = 4667
    #10;
    addra = 32'd149376;
    dina = {96'd0, 16'd30923, 16'd25008, 16'd2263, 16'd41245, 16'd49495, 16'd33530, 16'd842, 16'd6911, 16'd42457, 16'd34343}; // indx = 4668
    #10;
    addra = 32'd149408;
    dina = {96'd0, 16'd64998, 16'd48780, 16'd37857, 16'd35715, 16'd1877, 16'd1789, 16'd39115, 16'd19664, 16'd49835, 16'd15276}; // indx = 4669
    #10;
    addra = 32'd149440;
    dina = {96'd0, 16'd8319, 16'd33556, 16'd48847, 16'd41407, 16'd28496, 16'd23550, 16'd43847, 16'd48677, 16'd45187, 16'd50951}; // indx = 4670
    #10;
    addra = 32'd149472;
    dina = {96'd0, 16'd42203, 16'd10893, 16'd56555, 16'd29671, 16'd56825, 16'd65174, 16'd42669, 16'd35390, 16'd13416, 16'd57947}; // indx = 4671
    #10;
    addra = 32'd149504;
    dina = {96'd0, 16'd14492, 16'd16317, 16'd41694, 16'd46734, 16'd39652, 16'd17506, 16'd53723, 16'd12683, 16'd14469, 16'd60033}; // indx = 4672
    #10;
    addra = 32'd149536;
    dina = {96'd0, 16'd16592, 16'd34360, 16'd27836, 16'd25169, 16'd44050, 16'd9043, 16'd23723, 16'd16467, 16'd2834, 16'd15662}; // indx = 4673
    #10;
    addra = 32'd149568;
    dina = {96'd0, 16'd34458, 16'd46186, 16'd1015, 16'd25804, 16'd41212, 16'd2631, 16'd16004, 16'd10685, 16'd266, 16'd35722}; // indx = 4674
    #10;
    addra = 32'd149600;
    dina = {96'd0, 16'd37645, 16'd39948, 16'd55367, 16'd51754, 16'd8892, 16'd19868, 16'd4288, 16'd16191, 16'd48344, 16'd30946}; // indx = 4675
    #10;
    addra = 32'd149632;
    dina = {96'd0, 16'd27369, 16'd46723, 16'd59233, 16'd22855, 16'd34136, 16'd31376, 16'd24551, 16'd39049, 16'd15067, 16'd11061}; // indx = 4676
    #10;
    addra = 32'd149664;
    dina = {96'd0, 16'd51302, 16'd53636, 16'd35200, 16'd50353, 16'd6699, 16'd55034, 16'd32635, 16'd36511, 16'd8359, 16'd43834}; // indx = 4677
    #10;
    addra = 32'd149696;
    dina = {96'd0, 16'd41501, 16'd53762, 16'd10072, 16'd4291, 16'd61634, 16'd62818, 16'd29727, 16'd26895, 16'd45116, 16'd12250}; // indx = 4678
    #10;
    addra = 32'd149728;
    dina = {96'd0, 16'd11438, 16'd40708, 16'd17381, 16'd56610, 16'd58160, 16'd29329, 16'd46656, 16'd42156, 16'd4708, 16'd25437}; // indx = 4679
    #10;
    addra = 32'd149760;
    dina = {96'd0, 16'd34868, 16'd44217, 16'd17633, 16'd42344, 16'd50901, 16'd59264, 16'd25208, 16'd38480, 16'd40188, 16'd24559}; // indx = 4680
    #10;
    addra = 32'd149792;
    dina = {96'd0, 16'd50512, 16'd2669, 16'd43669, 16'd53685, 16'd34356, 16'd45284, 16'd16281, 16'd33459, 16'd16499, 16'd34923}; // indx = 4681
    #10;
    addra = 32'd149824;
    dina = {96'd0, 16'd19364, 16'd34718, 16'd56635, 16'd52288, 16'd57979, 16'd47227, 16'd18281, 16'd37019, 16'd58904, 16'd15764}; // indx = 4682
    #10;
    addra = 32'd149856;
    dina = {96'd0, 16'd39482, 16'd9316, 16'd2066, 16'd49905, 16'd47522, 16'd52148, 16'd10428, 16'd24438, 16'd3680, 16'd59405}; // indx = 4683
    #10;
    addra = 32'd149888;
    dina = {96'd0, 16'd6025, 16'd14975, 16'd22740, 16'd55728, 16'd42104, 16'd9352, 16'd41651, 16'd14880, 16'd26726, 16'd62918}; // indx = 4684
    #10;
    addra = 32'd149920;
    dina = {96'd0, 16'd56926, 16'd31575, 16'd4967, 16'd25936, 16'd42421, 16'd43508, 16'd44663, 16'd13891, 16'd53708, 16'd36752}; // indx = 4685
    #10;
    addra = 32'd149952;
    dina = {96'd0, 16'd56508, 16'd63300, 16'd50320, 16'd21493, 16'd25464, 16'd32459, 16'd18730, 16'd16158, 16'd41219, 16'd31230}; // indx = 4686
    #10;
    addra = 32'd149984;
    dina = {96'd0, 16'd11496, 16'd34826, 16'd62425, 16'd62324, 16'd7218, 16'd41244, 16'd51273, 16'd42719, 16'd48679, 16'd60293}; // indx = 4687
    #10;
    addra = 32'd150016;
    dina = {96'd0, 16'd42684, 16'd43083, 16'd58912, 16'd51532, 16'd21049, 16'd63570, 16'd27914, 16'd24248, 16'd59505, 16'd12228}; // indx = 4688
    #10;
    addra = 32'd150048;
    dina = {96'd0, 16'd30879, 16'd35363, 16'd49327, 16'd18048, 16'd65375, 16'd47935, 16'd24294, 16'd58176, 16'd19044, 16'd62589}; // indx = 4689
    #10;
    addra = 32'd150080;
    dina = {96'd0, 16'd61602, 16'd47378, 16'd58471, 16'd27244, 16'd58673, 16'd13389, 16'd11878, 16'd23419, 16'd10297, 16'd37657}; // indx = 4690
    #10;
    addra = 32'd150112;
    dina = {96'd0, 16'd1737, 16'd20262, 16'd7892, 16'd48587, 16'd52296, 16'd61661, 16'd62501, 16'd41084, 16'd57318, 16'd21915}; // indx = 4691
    #10;
    addra = 32'd150144;
    dina = {96'd0, 16'd59415, 16'd47477, 16'd23367, 16'd10405, 16'd17704, 16'd29139, 16'd60646, 16'd13099, 16'd62608, 16'd56934}; // indx = 4692
    #10;
    addra = 32'd150176;
    dina = {96'd0, 16'd13315, 16'd46954, 16'd5606, 16'd18213, 16'd19850, 16'd56404, 16'd45532, 16'd15759, 16'd10379, 16'd61049}; // indx = 4693
    #10;
    addra = 32'd150208;
    dina = {96'd0, 16'd64390, 16'd997, 16'd38746, 16'd29525, 16'd47502, 16'd22639, 16'd35198, 16'd16723, 16'd21963, 16'd21292}; // indx = 4694
    #10;
    addra = 32'd150240;
    dina = {96'd0, 16'd24789, 16'd34854, 16'd21663, 16'd27995, 16'd16290, 16'd9813, 16'd41275, 16'd19698, 16'd65197, 16'd5807}; // indx = 4695
    #10;
    addra = 32'd150272;
    dina = {96'd0, 16'd28352, 16'd42856, 16'd42255, 16'd51167, 16'd9644, 16'd59099, 16'd52995, 16'd55286, 16'd58030, 16'd38474}; // indx = 4696
    #10;
    addra = 32'd150304;
    dina = {96'd0, 16'd32747, 16'd38091, 16'd38682, 16'd38116, 16'd52754, 16'd60756, 16'd8160, 16'd15172, 16'd30951, 16'd53849}; // indx = 4697
    #10;
    addra = 32'd150336;
    dina = {96'd0, 16'd42188, 16'd10189, 16'd38751, 16'd33634, 16'd8557, 16'd62560, 16'd28695, 16'd34253, 16'd12374, 16'd23841}; // indx = 4698
    #10;
    addra = 32'd150368;
    dina = {96'd0, 16'd10565, 16'd14507, 16'd16123, 16'd19889, 16'd54454, 16'd29156, 16'd60131, 16'd37174, 16'd16315, 16'd43722}; // indx = 4699
    #10;
    addra = 32'd150400;
    dina = {96'd0, 16'd25228, 16'd50068, 16'd13191, 16'd58528, 16'd5494, 16'd43075, 16'd48071, 16'd20928, 16'd9044, 16'd6862}; // indx = 4700
    #10;
    addra = 32'd150432;
    dina = {96'd0, 16'd30895, 16'd42185, 16'd65343, 16'd50299, 16'd5408, 16'd62530, 16'd45057, 16'd125, 16'd21320, 16'd55785}; // indx = 4701
    #10;
    addra = 32'd150464;
    dina = {96'd0, 16'd57359, 16'd14028, 16'd32282, 16'd11568, 16'd50888, 16'd37391, 16'd8350, 16'd62394, 16'd60645, 16'd41792}; // indx = 4702
    #10;
    addra = 32'd150496;
    dina = {96'd0, 16'd63210, 16'd19989, 16'd62879, 16'd20890, 16'd4116, 16'd24088, 16'd60342, 16'd12784, 16'd34670, 16'd34246}; // indx = 4703
    #10;
    addra = 32'd150528;
    dina = {96'd0, 16'd14828, 16'd41431, 16'd16607, 16'd8087, 16'd14161, 16'd24406, 16'd31676, 16'd6084, 16'd44108, 16'd63061}; // indx = 4704
    #10;
    addra = 32'd150560;
    dina = {96'd0, 16'd52737, 16'd14892, 16'd37373, 16'd41976, 16'd38307, 16'd56214, 16'd64103, 16'd23557, 16'd17278, 16'd41983}; // indx = 4705
    #10;
    addra = 32'd150592;
    dina = {96'd0, 16'd3581, 16'd29826, 16'd13084, 16'd42445, 16'd45051, 16'd51712, 16'd61720, 16'd62781, 16'd1835, 16'd21104}; // indx = 4706
    #10;
    addra = 32'd150624;
    dina = {96'd0, 16'd12530, 16'd8904, 16'd61265, 16'd21691, 16'd16148, 16'd13778, 16'd12414, 16'd56861, 16'd55618, 16'd61610}; // indx = 4707
    #10;
    addra = 32'd150656;
    dina = {96'd0, 16'd64109, 16'd49772, 16'd37543, 16'd27600, 16'd33275, 16'd34823, 16'd55787, 16'd21098, 16'd33408, 16'd46797}; // indx = 4708
    #10;
    addra = 32'd150688;
    dina = {96'd0, 16'd5631, 16'd44504, 16'd22563, 16'd29939, 16'd30101, 16'd32781, 16'd37764, 16'd7839, 16'd64430, 16'd35055}; // indx = 4709
    #10;
    addra = 32'd150720;
    dina = {96'd0, 16'd47221, 16'd37495, 16'd10991, 16'd46122, 16'd13133, 16'd11637, 16'd29484, 16'd22824, 16'd1856, 16'd51507}; // indx = 4710
    #10;
    addra = 32'd150752;
    dina = {96'd0, 16'd48553, 16'd35508, 16'd42439, 16'd10803, 16'd7372, 16'd4195, 16'd56437, 16'd6086, 16'd12922, 16'd6796}; // indx = 4711
    #10;
    addra = 32'd150784;
    dina = {96'd0, 16'd1189, 16'd63379, 16'd6979, 16'd48374, 16'd5279, 16'd15669, 16'd9344, 16'd53306, 16'd30181, 16'd56828}; // indx = 4712
    #10;
    addra = 32'd150816;
    dina = {96'd0, 16'd26053, 16'd41471, 16'd24322, 16'd60566, 16'd64626, 16'd56054, 16'd14440, 16'd39691, 16'd63154, 16'd22057}; // indx = 4713
    #10;
    addra = 32'd150848;
    dina = {96'd0, 16'd48277, 16'd48347, 16'd6840, 16'd53160, 16'd54898, 16'd30033, 16'd10264, 16'd2699, 16'd27565, 16'd59271}; // indx = 4714
    #10;
    addra = 32'd150880;
    dina = {96'd0, 16'd9168, 16'd32323, 16'd64645, 16'd23051, 16'd14132, 16'd2501, 16'd49472, 16'd51107, 16'd11877, 16'd3410}; // indx = 4715
    #10;
    addra = 32'd150912;
    dina = {96'd0, 16'd9154, 16'd43219, 16'd39011, 16'd44119, 16'd14495, 16'd25032, 16'd11919, 16'd60486, 16'd39537, 16'd54514}; // indx = 4716
    #10;
    addra = 32'd150944;
    dina = {96'd0, 16'd41287, 16'd47960, 16'd27610, 16'd15270, 16'd11015, 16'd37461, 16'd51155, 16'd21741, 16'd14659, 16'd31767}; // indx = 4717
    #10;
    addra = 32'd150976;
    dina = {96'd0, 16'd40845, 16'd1872, 16'd42666, 16'd60730, 16'd10269, 16'd9045, 16'd4696, 16'd2176, 16'd39004, 16'd39602}; // indx = 4718
    #10;
    addra = 32'd151008;
    dina = {96'd0, 16'd2615, 16'd32128, 16'd31688, 16'd9666, 16'd11091, 16'd19420, 16'd638, 16'd61903, 16'd11995, 16'd18448}; // indx = 4719
    #10;
    addra = 32'd151040;
    dina = {96'd0, 16'd42010, 16'd39908, 16'd57767, 16'd49059, 16'd51139, 16'd19747, 16'd20706, 16'd1453, 16'd35707, 16'd26469}; // indx = 4720
    #10;
    addra = 32'd151072;
    dina = {96'd0, 16'd44785, 16'd29490, 16'd4474, 16'd20995, 16'd38350, 16'd52743, 16'd12651, 16'd58216, 16'd24676, 16'd29036}; // indx = 4721
    #10;
    addra = 32'd151104;
    dina = {96'd0, 16'd36959, 16'd60465, 16'd2430, 16'd21657, 16'd55782, 16'd46599, 16'd32413, 16'd30925, 16'd41658, 16'd52935}; // indx = 4722
    #10;
    addra = 32'd151136;
    dina = {96'd0, 16'd61069, 16'd11182, 16'd40953, 16'd36109, 16'd571, 16'd17626, 16'd40360, 16'd13960, 16'd217, 16'd13397}; // indx = 4723
    #10;
    addra = 32'd151168;
    dina = {96'd0, 16'd43237, 16'd38931, 16'd45081, 16'd30371, 16'd10467, 16'd36906, 16'd9925, 16'd59290, 16'd22624, 16'd18564}; // indx = 4724
    #10;
    addra = 32'd151200;
    dina = {96'd0, 16'd26731, 16'd19559, 16'd10944, 16'd57952, 16'd56480, 16'd29160, 16'd32554, 16'd7496, 16'd15428, 16'd43643}; // indx = 4725
    #10;
    addra = 32'd151232;
    dina = {96'd0, 16'd50463, 16'd2976, 16'd49722, 16'd40053, 16'd57978, 16'd37244, 16'd25626, 16'd3446, 16'd49714, 16'd60870}; // indx = 4726
    #10;
    addra = 32'd151264;
    dina = {96'd0, 16'd50557, 16'd3149, 16'd27688, 16'd60383, 16'd48502, 16'd24460, 16'd20185, 16'd46341, 16'd47344, 16'd65094}; // indx = 4727
    #10;
    addra = 32'd151296;
    dina = {96'd0, 16'd51172, 16'd16259, 16'd29274, 16'd26943, 16'd33827, 16'd49268, 16'd17907, 16'd9569, 16'd40405, 16'd38471}; // indx = 4728
    #10;
    addra = 32'd151328;
    dina = {96'd0, 16'd26958, 16'd37794, 16'd56386, 16'd21476, 16'd17117, 16'd59458, 16'd36000, 16'd2833, 16'd25935, 16'd11237}; // indx = 4729
    #10;
    addra = 32'd151360;
    dina = {96'd0, 16'd38899, 16'd30107, 16'd44774, 16'd59173, 16'd16255, 16'd34997, 16'd27299, 16'd42397, 16'd20211, 16'd863}; // indx = 4730
    #10;
    addra = 32'd151392;
    dina = {96'd0, 16'd584, 16'd59534, 16'd18737, 16'd8303, 16'd63374, 16'd6278, 16'd63751, 16'd17118, 16'd35808, 16'd21721}; // indx = 4731
    #10;
    addra = 32'd151424;
    dina = {96'd0, 16'd1169, 16'd27467, 16'd63789, 16'd22767, 16'd6834, 16'd50032, 16'd31515, 16'd5617, 16'd12875, 16'd54595}; // indx = 4732
    #10;
    addra = 32'd151456;
    dina = {96'd0, 16'd49481, 16'd31895, 16'd32654, 16'd6932, 16'd54471, 16'd43557, 16'd55536, 16'd4940, 16'd47460, 16'd20361}; // indx = 4733
    #10;
    addra = 32'd151488;
    dina = {96'd0, 16'd63515, 16'd47828, 16'd56069, 16'd63434, 16'd35071, 16'd16756, 16'd9468, 16'd48423, 16'd15167, 16'd35720}; // indx = 4734
    #10;
    addra = 32'd151520;
    dina = {96'd0, 16'd30836, 16'd55585, 16'd40373, 16'd62927, 16'd8465, 16'd5876, 16'd40244, 16'd27370, 16'd56357, 16'd3828}; // indx = 4735
    #10;
    addra = 32'd151552;
    dina = {96'd0, 16'd30171, 16'd28171, 16'd35441, 16'd48858, 16'd1402, 16'd23186, 16'd8472, 16'd19625, 16'd51802, 16'd45550}; // indx = 4736
    #10;
    addra = 32'd151584;
    dina = {96'd0, 16'd17496, 16'd61320, 16'd4847, 16'd8947, 16'd895, 16'd15659, 16'd32339, 16'd64777, 16'd19143, 16'd48416}; // indx = 4737
    #10;
    addra = 32'd151616;
    dina = {96'd0, 16'd16912, 16'd42915, 16'd21217, 16'd953, 16'd29968, 16'd18794, 16'd43754, 16'd39803, 16'd630, 16'd33635}; // indx = 4738
    #10;
    addra = 32'd151648;
    dina = {96'd0, 16'd24693, 16'd21214, 16'd24052, 16'd6365, 16'd31963, 16'd63721, 16'd23915, 16'd65231, 16'd6428, 16'd41258}; // indx = 4739
    #10;
    addra = 32'd151680;
    dina = {96'd0, 16'd16041, 16'd59674, 16'd46040, 16'd65146, 16'd28095, 16'd59669, 16'd38939, 16'd65030, 16'd54579, 16'd29087}; // indx = 4740
    #10;
    addra = 32'd151712;
    dina = {96'd0, 16'd23133, 16'd51082, 16'd63257, 16'd60677, 16'd20598, 16'd28278, 16'd17866, 16'd13011, 16'd65149, 16'd21649}; // indx = 4741
    #10;
    addra = 32'd151744;
    dina = {96'd0, 16'd23833, 16'd20935, 16'd27741, 16'd51434, 16'd1788, 16'd13680, 16'd50666, 16'd40718, 16'd48255, 16'd7248}; // indx = 4742
    #10;
    addra = 32'd151776;
    dina = {96'd0, 16'd33178, 16'd45261, 16'd27761, 16'd19980, 16'd18857, 16'd50720, 16'd8003, 16'd41828, 16'd55769, 16'd64690}; // indx = 4743
    #10;
    addra = 32'd151808;
    dina = {96'd0, 16'd38771, 16'd16944, 16'd65227, 16'd15881, 16'd8981, 16'd1549, 16'd47848, 16'd27103, 16'd31544, 16'd22550}; // indx = 4744
    #10;
    addra = 32'd151840;
    dina = {96'd0, 16'd20974, 16'd7881, 16'd12445, 16'd44399, 16'd39494, 16'd61203, 16'd42383, 16'd38820, 16'd26524, 16'd7818}; // indx = 4745
    #10;
    addra = 32'd151872;
    dina = {96'd0, 16'd61776, 16'd19397, 16'd65493, 16'd15646, 16'd56681, 16'd6345, 16'd53021, 16'd4812, 16'd1324, 16'd8173}; // indx = 4746
    #10;
    addra = 32'd151904;
    dina = {96'd0, 16'd36381, 16'd54278, 16'd12648, 16'd43695, 16'd871, 16'd23877, 16'd26120, 16'd41869, 16'd29195, 16'd36268}; // indx = 4747
    #10;
    addra = 32'd151936;
    dina = {96'd0, 16'd44990, 16'd5384, 16'd11040, 16'd8664, 16'd43806, 16'd7671, 16'd35798, 16'd15686, 16'd20861, 16'd7013}; // indx = 4748
    #10;
    addra = 32'd151968;
    dina = {96'd0, 16'd36436, 16'd17123, 16'd4507, 16'd41453, 16'd14066, 16'd14119, 16'd28823, 16'd7009, 16'd2699, 16'd36365}; // indx = 4749
    #10;
    addra = 32'd152000;
    dina = {96'd0, 16'd1387, 16'd32396, 16'd39334, 16'd65425, 16'd30482, 16'd62047, 16'd19712, 16'd51193, 16'd1326, 16'd39129}; // indx = 4750
    #10;
    addra = 32'd152032;
    dina = {96'd0, 16'd32860, 16'd13735, 16'd26728, 16'd9531, 16'd33960, 16'd43192, 16'd43206, 16'd42786, 16'd37920, 16'd40702}; // indx = 4751
    #10;
    addra = 32'd152064;
    dina = {96'd0, 16'd12441, 16'd31078, 16'd18853, 16'd25136, 16'd43123, 16'd40666, 16'd49976, 16'd15077, 16'd51474, 16'd230}; // indx = 4752
    #10;
    addra = 32'd152096;
    dina = {96'd0, 16'd45299, 16'd28119, 16'd9969, 16'd15294, 16'd35059, 16'd38525, 16'd55277, 16'd37882, 16'd40456, 16'd18161}; // indx = 4753
    #10;
    addra = 32'd152128;
    dina = {96'd0, 16'd20014, 16'd11470, 16'd61189, 16'd15493, 16'd337, 16'd17947, 16'd39697, 16'd11434, 16'd11331, 16'd64552}; // indx = 4754
    #10;
    addra = 32'd152160;
    dina = {96'd0, 16'd60993, 16'd27826, 16'd3153, 16'd48536, 16'd47486, 16'd19227, 16'd4649, 16'd57972, 16'd3862, 16'd60148}; // indx = 4755
    #10;
    addra = 32'd152192;
    dina = {96'd0, 16'd23620, 16'd24553, 16'd35059, 16'd54999, 16'd11365, 16'd61841, 16'd8025, 16'd54788, 16'd34497, 16'd31470}; // indx = 4756
    #10;
    addra = 32'd152224;
    dina = {96'd0, 16'd15455, 16'd5648, 16'd5599, 16'd51073, 16'd41158, 16'd15435, 16'd30144, 16'd54179, 16'd43831, 16'd6730}; // indx = 4757
    #10;
    addra = 32'd152256;
    dina = {96'd0, 16'd49570, 16'd25016, 16'd41769, 16'd39983, 16'd8741, 16'd35896, 16'd13795, 16'd37420, 16'd14684, 16'd25605}; // indx = 4758
    #10;
    addra = 32'd152288;
    dina = {96'd0, 16'd52864, 16'd52287, 16'd37488, 16'd61663, 16'd63834, 16'd15064, 16'd18068, 16'd8999, 16'd52393, 16'd60936}; // indx = 4759
    #10;
    addra = 32'd152320;
    dina = {96'd0, 16'd16368, 16'd45492, 16'd28204, 16'd34744, 16'd13517, 16'd64040, 16'd58181, 16'd40456, 16'd53867, 16'd5156}; // indx = 4760
    #10;
    addra = 32'd152352;
    dina = {96'd0, 16'd5273, 16'd18990, 16'd47130, 16'd63087, 16'd44096, 16'd42737, 16'd55368, 16'd42598, 16'd35077, 16'd45736}; // indx = 4761
    #10;
    addra = 32'd152384;
    dina = {96'd0, 16'd31190, 16'd52182, 16'd32828, 16'd5703, 16'd2072, 16'd45621, 16'd60391, 16'd14438, 16'd61348, 16'd17011}; // indx = 4762
    #10;
    addra = 32'd152416;
    dina = {96'd0, 16'd9695, 16'd41452, 16'd21051, 16'd7400, 16'd36650, 16'd45396, 16'd47242, 16'd56025, 16'd40438, 16'd38422}; // indx = 4763
    #10;
    addra = 32'd152448;
    dina = {96'd0, 16'd49564, 16'd32407, 16'd36090, 16'd4162, 16'd44148, 16'd5058, 16'd33777, 16'd41790, 16'd21749, 16'd18645}; // indx = 4764
    #10;
    addra = 32'd152480;
    dina = {96'd0, 16'd40557, 16'd63467, 16'd13171, 16'd52023, 16'd37461, 16'd39334, 16'd47893, 16'd47326, 16'd16812, 16'd33592}; // indx = 4765
    #10;
    addra = 32'd152512;
    dina = {96'd0, 16'd62822, 16'd15306, 16'd21406, 16'd11363, 16'd58179, 16'd145, 16'd1429, 16'd7748, 16'd50760, 16'd42338}; // indx = 4766
    #10;
    addra = 32'd152544;
    dina = {96'd0, 16'd56989, 16'd40058, 16'd43102, 16'd24940, 16'd58949, 16'd10303, 16'd59410, 16'd52313, 16'd4146, 16'd36921}; // indx = 4767
    #10;
    addra = 32'd152576;
    dina = {96'd0, 16'd27350, 16'd36967, 16'd43387, 16'd43232, 16'd53040, 16'd23468, 16'd20006, 16'd64732, 16'd59980, 16'd50419}; // indx = 4768
    #10;
    addra = 32'd152608;
    dina = {96'd0, 16'd17383, 16'd34684, 16'd38717, 16'd4275, 16'd16480, 16'd10547, 16'd35097, 16'd61010, 16'd58198, 16'd63184}; // indx = 4769
    #10;
    addra = 32'd152640;
    dina = {96'd0, 16'd50701, 16'd62615, 16'd15069, 16'd54360, 16'd29996, 16'd3976, 16'd18497, 16'd61947, 16'd62379, 16'd37170}; // indx = 4770
    #10;
    addra = 32'd152672;
    dina = {96'd0, 16'd59914, 16'd1931, 16'd24714, 16'd33273, 16'd20133, 16'd57921, 16'd17222, 16'd55907, 16'd3551, 16'd59393}; // indx = 4771
    #10;
    addra = 32'd152704;
    dina = {96'd0, 16'd54779, 16'd41398, 16'd42913, 16'd27821, 16'd39313, 16'd16983, 16'd26251, 16'd44790, 16'd31631, 16'd27567}; // indx = 4772
    #10;
    addra = 32'd152736;
    dina = {96'd0, 16'd43454, 16'd29016, 16'd4458, 16'd19355, 16'd38506, 16'd35071, 16'd25221, 16'd36998, 16'd56613, 16'd40334}; // indx = 4773
    #10;
    addra = 32'd152768;
    dina = {96'd0, 16'd53340, 16'd24598, 16'd28946, 16'd52197, 16'd8367, 16'd14225, 16'd35722, 16'd24318, 16'd26208, 16'd61601}; // indx = 4774
    #10;
    addra = 32'd152800;
    dina = {96'd0, 16'd52502, 16'd49492, 16'd19502, 16'd52841, 16'd16846, 16'd44093, 16'd54733, 16'd65182, 16'd62524, 16'd59050}; // indx = 4775
    #10;
    addra = 32'd152832;
    dina = {96'd0, 16'd65487, 16'd23019, 16'd62641, 16'd28048, 16'd45267, 16'd61130, 16'd56994, 16'd36492, 16'd60267, 16'd38980}; // indx = 4776
    #10;
    addra = 32'd152864;
    dina = {96'd0, 16'd28899, 16'd27076, 16'd37881, 16'd55892, 16'd17960, 16'd39256, 16'd33625, 16'd61158, 16'd1402, 16'd36926}; // indx = 4777
    #10;
    addra = 32'd152896;
    dina = {96'd0, 16'd26942, 16'd58003, 16'd32449, 16'd22189, 16'd11261, 16'd28285, 16'd18952, 16'd26078, 16'd22968, 16'd49703}; // indx = 4778
    #10;
    addra = 32'd152928;
    dina = {96'd0, 16'd20447, 16'd56146, 16'd53906, 16'd8787, 16'd14653, 16'd6149, 16'd36031, 16'd18891, 16'd13282, 16'd29710}; // indx = 4779
    #10;
    addra = 32'd152960;
    dina = {96'd0, 16'd48696, 16'd17054, 16'd34946, 16'd2904, 16'd54296, 16'd50859, 16'd7042, 16'd40553, 16'd15653, 16'd5238}; // indx = 4780
    #10;
    addra = 32'd152992;
    dina = {96'd0, 16'd43862, 16'd14815, 16'd33061, 16'd45135, 16'd59592, 16'd28878, 16'd36963, 16'd13689, 16'd36784, 16'd29554}; // indx = 4781
    #10;
    addra = 32'd153024;
    dina = {96'd0, 16'd45057, 16'd57394, 16'd22372, 16'd44975, 16'd56699, 16'd24717, 16'd11860, 16'd54251, 16'd14731, 16'd40029}; // indx = 4782
    #10;
    addra = 32'd153056;
    dina = {96'd0, 16'd34844, 16'd44229, 16'd20404, 16'd56586, 16'd17496, 16'd46044, 16'd34587, 16'd25153, 16'd50198, 16'd47519}; // indx = 4783
    #10;
    addra = 32'd153088;
    dina = {96'd0, 16'd52936, 16'd19845, 16'd4947, 16'd58068, 16'd23386, 16'd4826, 16'd39595, 16'd19412, 16'd55799, 16'd29898}; // indx = 4784
    #10;
    addra = 32'd153120;
    dina = {96'd0, 16'd16024, 16'd51320, 16'd27225, 16'd49643, 16'd12374, 16'd13167, 16'd58964, 16'd15868, 16'd57812, 16'd35265}; // indx = 4785
    #10;
    addra = 32'd153152;
    dina = {96'd0, 16'd37009, 16'd45632, 16'd53285, 16'd39439, 16'd51245, 16'd2034, 16'd34878, 16'd17444, 16'd10771, 16'd20729}; // indx = 4786
    #10;
    addra = 32'd153184;
    dina = {96'd0, 16'd19246, 16'd54025, 16'd15052, 16'd31037, 16'd56195, 16'd24086, 16'd53907, 16'd18348, 16'd58542, 16'd5577}; // indx = 4787
    #10;
    addra = 32'd153216;
    dina = {96'd0, 16'd3619, 16'd39349, 16'd20462, 16'd17686, 16'd6087, 16'd35840, 16'd23701, 16'd33690, 16'd27634, 16'd52341}; // indx = 4788
    #10;
    addra = 32'd153248;
    dina = {96'd0, 16'd4198, 16'd36867, 16'd26203, 16'd42046, 16'd48348, 16'd45014, 16'd53559, 16'd58733, 16'd44092, 16'd18453}; // indx = 4789
    #10;
    addra = 32'd153280;
    dina = {96'd0, 16'd28352, 16'd48330, 16'd52032, 16'd10058, 16'd44578, 16'd12510, 16'd28752, 16'd62652, 16'd33486, 16'd62984}; // indx = 4790
    #10;
    addra = 32'd153312;
    dina = {96'd0, 16'd64310, 16'd22518, 16'd10099, 16'd28729, 16'd20435, 16'd19927, 16'd54568, 16'd8684, 16'd40823, 16'd19478}; // indx = 4791
    #10;
    addra = 32'd153344;
    dina = {96'd0, 16'd43615, 16'd39035, 16'd64281, 16'd15422, 16'd27537, 16'd2084, 16'd41779, 16'd31359, 16'd9301, 16'd16057}; // indx = 4792
    #10;
    addra = 32'd153376;
    dina = {96'd0, 16'd31305, 16'd55616, 16'd13599, 16'd17865, 16'd41853, 16'd23111, 16'd24802, 16'd49688, 16'd4472, 16'd29993}; // indx = 4793
    #10;
    addra = 32'd153408;
    dina = {96'd0, 16'd7307, 16'd4134, 16'd33687, 16'd45517, 16'd20827, 16'd58648, 16'd11762, 16'd37778, 16'd37454, 16'd51227}; // indx = 4794
    #10;
    addra = 32'd153440;
    dina = {96'd0, 16'd39924, 16'd732, 16'd45692, 16'd57365, 16'd6876, 16'd33803, 16'd12391, 16'd30567, 16'd18515, 16'd6595}; // indx = 4795
    #10;
    addra = 32'd153472;
    dina = {96'd0, 16'd7009, 16'd61245, 16'd62146, 16'd9599, 16'd28281, 16'd60565, 16'd24147, 16'd41381, 16'd53593, 16'd18875}; // indx = 4796
    #10;
    addra = 32'd153504;
    dina = {96'd0, 16'd18326, 16'd16954, 16'd3765, 16'd45911, 16'd9035, 16'd39385, 16'd59583, 16'd32959, 16'd65424, 16'd48795}; // indx = 4797
    #10;
    addra = 32'd153536;
    dina = {96'd0, 16'd6177, 16'd23800, 16'd15389, 16'd22107, 16'd60355, 16'd27840, 16'd28853, 16'd32161, 16'd32422, 16'd11796}; // indx = 4798
    #10;
    addra = 32'd153568;
    dina = {96'd0, 16'd13459, 16'd36931, 16'd31769, 16'd33780, 16'd15966, 16'd2195, 16'd54739, 16'd13450, 16'd32037, 16'd49101}; // indx = 4799
    #10;
    addra = 32'd153600;
    dina = {96'd0, 16'd41341, 16'd34860, 16'd11845, 16'd30603, 16'd58006, 16'd5827, 16'd27942, 16'd21979, 16'd26869, 16'd41526}; // indx = 4800
    #10;
    addra = 32'd153632;
    dina = {96'd0, 16'd26983, 16'd27788, 16'd12274, 16'd44463, 16'd42853, 16'd31374, 16'd10857, 16'd10063, 16'd65055, 16'd56079}; // indx = 4801
    #10;
    addra = 32'd153664;
    dina = {96'd0, 16'd6932, 16'd32660, 16'd8086, 16'd65320, 16'd29958, 16'd4217, 16'd5995, 16'd50961, 16'd22564, 16'd62803}; // indx = 4802
    #10;
    addra = 32'd153696;
    dina = {96'd0, 16'd36200, 16'd41609, 16'd35177, 16'd2005, 16'd23947, 16'd31783, 16'd32669, 16'd38804, 16'd47425, 16'd58734}; // indx = 4803
    #10;
    addra = 32'd153728;
    dina = {96'd0, 16'd18905, 16'd59745, 16'd34625, 16'd57437, 16'd53009, 16'd8001, 16'd36265, 16'd65516, 16'd49496, 16'd51431}; // indx = 4804
    #10;
    addra = 32'd153760;
    dina = {96'd0, 16'd27914, 16'd50719, 16'd9442, 16'd12469, 16'd14228, 16'd17634, 16'd17705, 16'd26598, 16'd54337, 16'd40729}; // indx = 4805
    #10;
    addra = 32'd153792;
    dina = {96'd0, 16'd13713, 16'd17216, 16'd16584, 16'd29726, 16'd48257, 16'd9591, 16'd64548, 16'd107, 16'd6835, 16'd28682}; // indx = 4806
    #10;
    addra = 32'd153824;
    dina = {96'd0, 16'd18349, 16'd5196, 16'd58510, 16'd52859, 16'd32449, 16'd42478, 16'd12980, 16'd16079, 16'd47246, 16'd41862}; // indx = 4807
    #10;
    addra = 32'd153856;
    dina = {96'd0, 16'd48121, 16'd65380, 16'd36403, 16'd34888, 16'd34726, 16'd45871, 16'd60097, 16'd59831, 16'd47684, 16'd1240}; // indx = 4808
    #10;
    addra = 32'd153888;
    dina = {96'd0, 16'd19808, 16'd22523, 16'd43462, 16'd11946, 16'd50828, 16'd22688, 16'd39036, 16'd53976, 16'd17461, 16'd36877}; // indx = 4809
    #10;
    addra = 32'd153920;
    dina = {96'd0, 16'd34879, 16'd1116, 16'd36636, 16'd9865, 16'd51555, 16'd47520, 16'd24446, 16'd31194, 16'd30327, 16'd24075}; // indx = 4810
    #10;
    addra = 32'd153952;
    dina = {96'd0, 16'd4539, 16'd63817, 16'd57253, 16'd21953, 16'd31125, 16'd11320, 16'd65064, 16'd62909, 16'd19256, 16'd23430}; // indx = 4811
    #10;
    addra = 32'd153984;
    dina = {96'd0, 16'd18546, 16'd10376, 16'd7950, 16'd13555, 16'd28741, 16'd7849, 16'd36983, 16'd56675, 16'd34693, 16'd31171}; // indx = 4812
    #10;
    addra = 32'd154016;
    dina = {96'd0, 16'd9491, 16'd63040, 16'd55265, 16'd24735, 16'd40819, 16'd55268, 16'd65377, 16'd48319, 16'd38221, 16'd58785}; // indx = 4813
    #10;
    addra = 32'd154048;
    dina = {96'd0, 16'd38948, 16'd16833, 16'd62386, 16'd9561, 16'd9581, 16'd46813, 16'd30525, 16'd17684, 16'd30325, 16'd7961}; // indx = 4814
    #10;
    addra = 32'd154080;
    dina = {96'd0, 16'd64254, 16'd8382, 16'd27467, 16'd59191, 16'd28772, 16'd21916, 16'd22134, 16'd46326, 16'd996, 16'd19554}; // indx = 4815
    #10;
    addra = 32'd154112;
    dina = {96'd0, 16'd929, 16'd427, 16'd31028, 16'd7903, 16'd23430, 16'd28394, 16'd9755, 16'd33845, 16'd9171, 16'd23721}; // indx = 4816
    #10;
    addra = 32'd154144;
    dina = {96'd0, 16'd10698, 16'd24219, 16'd8084, 16'd46427, 16'd26342, 16'd28524, 16'd27320, 16'd64717, 16'd43138, 16'd36995}; // indx = 4817
    #10;
    addra = 32'd154176;
    dina = {96'd0, 16'd49751, 16'd40457, 16'd49990, 16'd17275, 16'd38700, 16'd46890, 16'd22660, 16'd51786, 16'd37480, 16'd32609}; // indx = 4818
    #10;
    addra = 32'd154208;
    dina = {96'd0, 16'd18993, 16'd44136, 16'd11237, 16'd60884, 16'd23321, 16'd18503, 16'd50005, 16'd985, 16'd53598, 16'd2823}; // indx = 4819
    #10;
    addra = 32'd154240;
    dina = {96'd0, 16'd24367, 16'd60584, 16'd16766, 16'd52931, 16'd42145, 16'd22243, 16'd21167, 16'd53873, 16'd30544, 16'd20338}; // indx = 4820
    #10;
    addra = 32'd154272;
    dina = {96'd0, 16'd62995, 16'd49023, 16'd22239, 16'd49818, 16'd39370, 16'd3772, 16'd2936, 16'd37687, 16'd23397, 16'd24892}; // indx = 4821
    #10;
    addra = 32'd154304;
    dina = {96'd0, 16'd56917, 16'd33991, 16'd31261, 16'd1893, 16'd51439, 16'd65056, 16'd41311, 16'd31850, 16'd17275, 16'd30057}; // indx = 4822
    #10;
    addra = 32'd154336;
    dina = {96'd0, 16'd47739, 16'd48735, 16'd38686, 16'd44189, 16'd36103, 16'd24247, 16'd14809, 16'd40731, 16'd48673, 16'd25200}; // indx = 4823
    #10;
    addra = 32'd154368;
    dina = {96'd0, 16'd42134, 16'd18400, 16'd39053, 16'd14337, 16'd32688, 16'd21207, 16'd40768, 16'd35386, 16'd2087, 16'd63606}; // indx = 4824
    #10;
    addra = 32'd154400;
    dina = {96'd0, 16'd19057, 16'd3731, 16'd41950, 16'd3221, 16'd30191, 16'd6083, 16'd55636, 16'd5736, 16'd26138, 16'd57920}; // indx = 4825
    #10;
    addra = 32'd154432;
    dina = {96'd0, 16'd64559, 16'd8961, 16'd18535, 16'd52889, 16'd21544, 16'd22864, 16'd16139, 16'd53984, 16'd18176, 16'd11611}; // indx = 4826
    #10;
    addra = 32'd154464;
    dina = {96'd0, 16'd5369, 16'd64260, 16'd1690, 16'd28488, 16'd9778, 16'd56876, 16'd32955, 16'd59799, 16'd10845, 16'd922}; // indx = 4827
    #10;
    addra = 32'd154496;
    dina = {96'd0, 16'd53860, 16'd49321, 16'd31298, 16'd562, 16'd62869, 16'd5455, 16'd60969, 16'd7577, 16'd28784, 16'd53992}; // indx = 4828
    #10;
    addra = 32'd154528;
    dina = {96'd0, 16'd6252, 16'd45200, 16'd43321, 16'd59469, 16'd44059, 16'd49429, 16'd21768, 16'd1461, 16'd36190, 16'd13583}; // indx = 4829
    #10;
    addra = 32'd154560;
    dina = {96'd0, 16'd29941, 16'd32488, 16'd54877, 16'd29868, 16'd23403, 16'd21880, 16'd63485, 16'd29636, 16'd27202, 16'd38671}; // indx = 4830
    #10;
    addra = 32'd154592;
    dina = {96'd0, 16'd64314, 16'd2589, 16'd14806, 16'd25979, 16'd45427, 16'd29536, 16'd51205, 16'd7560, 16'd34018, 16'd20591}; // indx = 4831
    #10;
    addra = 32'd154624;
    dina = {96'd0, 16'd37743, 16'd12573, 16'd63011, 16'd52114, 16'd15891, 16'd18830, 16'd37942, 16'd21949, 16'd44172, 16'd34127}; // indx = 4832
    #10;
    addra = 32'd154656;
    dina = {96'd0, 16'd22144, 16'd54501, 16'd51142, 16'd21317, 16'd7653, 16'd11907, 16'd4839, 16'd17247, 16'd54630, 16'd24586}; // indx = 4833
    #10;
    addra = 32'd154688;
    dina = {96'd0, 16'd30110, 16'd32253, 16'd37205, 16'd58942, 16'd39128, 16'd43521, 16'd35591, 16'd602, 16'd9956, 16'd48441}; // indx = 4834
    #10;
    addra = 32'd154720;
    dina = {96'd0, 16'd22991, 16'd37494, 16'd31198, 16'd4078, 16'd36729, 16'd45478, 16'd41789, 16'd23931, 16'd48682, 16'd4114}; // indx = 4835
    #10;
    addra = 32'd154752;
    dina = {96'd0, 16'd9018, 16'd30600, 16'd62074, 16'd35793, 16'd11783, 16'd61884, 16'd57567, 16'd48457, 16'd49426, 16'd23285}; // indx = 4836
    #10;
    addra = 32'd154784;
    dina = {96'd0, 16'd25880, 16'd24699, 16'd49410, 16'd58524, 16'd42265, 16'd20458, 16'd54826, 16'd27576, 16'd18816, 16'd55829}; // indx = 4837
    #10;
    addra = 32'd154816;
    dina = {96'd0, 16'd39073, 16'd29765, 16'd31446, 16'd21506, 16'd36078, 16'd28276, 16'd59450, 16'd50613, 16'd47624, 16'd51374}; // indx = 4838
    #10;
    addra = 32'd154848;
    dina = {96'd0, 16'd48036, 16'd54024, 16'd63967, 16'd63662, 16'd50277, 16'd39151, 16'd64396, 16'd19833, 16'd23090, 16'd58565}; // indx = 4839
    #10;
    addra = 32'd154880;
    dina = {96'd0, 16'd29016, 16'd21762, 16'd55331, 16'd17530, 16'd55774, 16'd24257, 16'd31747, 16'd34310, 16'd40834, 16'd17596}; // indx = 4840
    #10;
    addra = 32'd154912;
    dina = {96'd0, 16'd48146, 16'd44313, 16'd29329, 16'd47197, 16'd3645, 16'd5146, 16'd56335, 16'd17595, 16'd37978, 16'd623}; // indx = 4841
    #10;
    addra = 32'd154944;
    dina = {96'd0, 16'd55222, 16'd54756, 16'd36397, 16'd47264, 16'd60910, 16'd16619, 16'd60987, 16'd82, 16'd52120, 16'd11080}; // indx = 4842
    #10;
    addra = 32'd154976;
    dina = {96'd0, 16'd45528, 16'd31981, 16'd59026, 16'd18491, 16'd56797, 16'd11131, 16'd38081, 16'd49440, 16'd34533, 16'd49640}; // indx = 4843
    #10;
    addra = 32'd155008;
    dina = {96'd0, 16'd42671, 16'd30871, 16'd64462, 16'd42082, 16'd12858, 16'd9987, 16'd38783, 16'd42244, 16'd63030, 16'd9880}; // indx = 4844
    #10;
    addra = 32'd155040;
    dina = {96'd0, 16'd9529, 16'd11162, 16'd54567, 16'd17308, 16'd45233, 16'd19394, 16'd6454, 16'd470, 16'd7211, 16'd42531}; // indx = 4845
    #10;
    addra = 32'd155072;
    dina = {96'd0, 16'd63089, 16'd20941, 16'd29964, 16'd19761, 16'd51834, 16'd33712, 16'd48697, 16'd62938, 16'd58445, 16'd33525}; // indx = 4846
    #10;
    addra = 32'd155104;
    dina = {96'd0, 16'd62522, 16'd44677, 16'd6566, 16'd60402, 16'd40500, 16'd12179, 16'd5824, 16'd35115, 16'd31051, 16'd5003}; // indx = 4847
    #10;
    addra = 32'd155136;
    dina = {96'd0, 16'd46803, 16'd16034, 16'd623, 16'd31407, 16'd16818, 16'd63501, 16'd4492, 16'd43509, 16'd22616, 16'd59661}; // indx = 4848
    #10;
    addra = 32'd155168;
    dina = {96'd0, 16'd27711, 16'd21833, 16'd2772, 16'd41659, 16'd26798, 16'd12541, 16'd20697, 16'd60959, 16'd58731, 16'd39602}; // indx = 4849
    #10;
    addra = 32'd155200;
    dina = {96'd0, 16'd9865, 16'd22349, 16'd24004, 16'd27097, 16'd15890, 16'd26111, 16'd47636, 16'd57206, 16'd51813, 16'd45730}; // indx = 4850
    #10;
    addra = 32'd155232;
    dina = {96'd0, 16'd31987, 16'd60881, 16'd26615, 16'd1710, 16'd28541, 16'd31621, 16'd36200, 16'd40338, 16'd18590, 16'd60015}; // indx = 4851
    #10;
    addra = 32'd155264;
    dina = {96'd0, 16'd43757, 16'd23049, 16'd50909, 16'd11957, 16'd61202, 16'd2314, 16'd41475, 16'd59158, 16'd40358, 16'd57173}; // indx = 4852
    #10;
    addra = 32'd155296;
    dina = {96'd0, 16'd60263, 16'd33144, 16'd2125, 16'd64554, 16'd25117, 16'd43613, 16'd23511, 16'd25453, 16'd12147, 16'd7805}; // indx = 4853
    #10;
    addra = 32'd155328;
    dina = {96'd0, 16'd43587, 16'd47662, 16'd27360, 16'd3019, 16'd43943, 16'd45387, 16'd63591, 16'd51056, 16'd50168, 16'd32645}; // indx = 4854
    #10;
    addra = 32'd155360;
    dina = {96'd0, 16'd57933, 16'd14481, 16'd21641, 16'd29497, 16'd29190, 16'd13010, 16'd34859, 16'd65398, 16'd40236, 16'd36057}; // indx = 4855
    #10;
    addra = 32'd155392;
    dina = {96'd0, 16'd64992, 16'd43626, 16'd62378, 16'd45761, 16'd49891, 16'd5608, 16'd41751, 16'd17620, 16'd18872, 16'd17781}; // indx = 4856
    #10;
    addra = 32'd155424;
    dina = {96'd0, 16'd44282, 16'd43494, 16'd30056, 16'd35978, 16'd33652, 16'd6490, 16'd24706, 16'd6115, 16'd24754, 16'd55926}; // indx = 4857
    #10;
    addra = 32'd155456;
    dina = {96'd0, 16'd899, 16'd54774, 16'd43510, 16'd13384, 16'd62400, 16'd7210, 16'd23609, 16'd8376, 16'd52587, 16'd59189}; // indx = 4858
    #10;
    addra = 32'd155488;
    dina = {96'd0, 16'd45137, 16'd39560, 16'd23210, 16'd30199, 16'd19324, 16'd51517, 16'd20214, 16'd55655, 16'd17261, 16'd20611}; // indx = 4859
    #10;
    addra = 32'd155520;
    dina = {96'd0, 16'd36867, 16'd49556, 16'd15630, 16'd11110, 16'd25878, 16'd2426, 16'd64919, 16'd50835, 16'd46020, 16'd14833}; // indx = 4860
    #10;
    addra = 32'd155552;
    dina = {96'd0, 16'd27881, 16'd3297, 16'd20038, 16'd44977, 16'd33210, 16'd3934, 16'd52253, 16'd44577, 16'd31090, 16'd30989}; // indx = 4861
    #10;
    addra = 32'd155584;
    dina = {96'd0, 16'd28782, 16'd15214, 16'd36923, 16'd61369, 16'd25266, 16'd37921, 16'd54948, 16'd41251, 16'd49291, 16'd42830}; // indx = 4862
    #10;
    addra = 32'd155616;
    dina = {96'd0, 16'd19524, 16'd30287, 16'd29264, 16'd13859, 16'd14626, 16'd56334, 16'd48798, 16'd57820, 16'd54152, 16'd62236}; // indx = 4863
    #10;
    addra = 32'd155648;
    dina = {96'd0, 16'd57039, 16'd38764, 16'd48224, 16'd37861, 16'd21737, 16'd63244, 16'd64354, 16'd4344, 16'd36044, 16'd16140}; // indx = 4864
    #10;
    addra = 32'd155680;
    dina = {96'd0, 16'd40633, 16'd2226, 16'd15424, 16'd18113, 16'd41050, 16'd43008, 16'd57801, 16'd30846, 16'd47975, 16'd9411}; // indx = 4865
    #10;
    addra = 32'd155712;
    dina = {96'd0, 16'd35098, 16'd57712, 16'd21080, 16'd52144, 16'd56893, 16'd10274, 16'd8890, 16'd63345, 16'd16860, 16'd16346}; // indx = 4866
    #10;
    addra = 32'd155744;
    dina = {96'd0, 16'd25456, 16'd37823, 16'd29516, 16'd50241, 16'd45698, 16'd51822, 16'd10449, 16'd7991, 16'd49337, 16'd49538}; // indx = 4867
    #10;
    addra = 32'd155776;
    dina = {96'd0, 16'd39344, 16'd62039, 16'd45631, 16'd677, 16'd27065, 16'd8284, 16'd26737, 16'd58679, 16'd26620, 16'd63646}; // indx = 4868
    #10;
    addra = 32'd155808;
    dina = {96'd0, 16'd17294, 16'd39707, 16'd53456, 16'd20720, 16'd47232, 16'd37734, 16'd38045, 16'd18734, 16'd14431, 16'd20588}; // indx = 4869
    #10;
    addra = 32'd155840;
    dina = {96'd0, 16'd20785, 16'd58263, 16'd659, 16'd63951, 16'd21708, 16'd8149, 16'd29596, 16'd40273, 16'd10401, 16'd5053}; // indx = 4870
    #10;
    addra = 32'd155872;
    dina = {96'd0, 16'd31025, 16'd38812, 16'd57334, 16'd24997, 16'd55833, 16'd32993, 16'd54052, 16'd23999, 16'd15205, 16'd18219}; // indx = 4871
    #10;
    addra = 32'd155904;
    dina = {96'd0, 16'd59307, 16'd47169, 16'd38643, 16'd40750, 16'd63077, 16'd19709, 16'd50219, 16'd60299, 16'd61843, 16'd61545}; // indx = 4872
    #10;
    addra = 32'd155936;
    dina = {96'd0, 16'd34649, 16'd6975, 16'd34028, 16'd38178, 16'd28540, 16'd55663, 16'd55884, 16'd4399, 16'd32118, 16'd63120}; // indx = 4873
    #10;
    addra = 32'd155968;
    dina = {96'd0, 16'd20900, 16'd54125, 16'd56302, 16'd56895, 16'd32872, 16'd45383, 16'd17092, 16'd524, 16'd26395, 16'd7232}; // indx = 4874
    #10;
    addra = 32'd156000;
    dina = {96'd0, 16'd35590, 16'd14725, 16'd19609, 16'd43012, 16'd54628, 16'd27342, 16'd17047, 16'd62320, 16'd14175, 16'd8767}; // indx = 4875
    #10;
    addra = 32'd156032;
    dina = {96'd0, 16'd33089, 16'd35869, 16'd61101, 16'd46030, 16'd44898, 16'd21162, 16'd21066, 16'd50278, 16'd29701, 16'd12334}; // indx = 4876
    #10;
    addra = 32'd156064;
    dina = {96'd0, 16'd42901, 16'd22259, 16'd43948, 16'd48741, 16'd37843, 16'd39601, 16'd17968, 16'd16770, 16'd56832, 16'd64294}; // indx = 4877
    #10;
    addra = 32'd156096;
    dina = {96'd0, 16'd11158, 16'd40595, 16'd19596, 16'd8850, 16'd41449, 16'd42696, 16'd11662, 16'd27751, 16'd37937, 16'd27518}; // indx = 4878
    #10;
    addra = 32'd156128;
    dina = {96'd0, 16'd54269, 16'd58983, 16'd7837, 16'd40268, 16'd47869, 16'd14467, 16'd53753, 16'd21711, 16'd40343, 16'd22038}; // indx = 4879
    #10;
    addra = 32'd156160;
    dina = {96'd0, 16'd31052, 16'd47852, 16'd15996, 16'd40623, 16'd31655, 16'd17558, 16'd13876, 16'd42699, 16'd4742, 16'd44562}; // indx = 4880
    #10;
    addra = 32'd156192;
    dina = {96'd0, 16'd25645, 16'd15063, 16'd27487, 16'd53667, 16'd17298, 16'd59284, 16'd1402, 16'd25522, 16'd59262, 16'd7623}; // indx = 4881
    #10;
    addra = 32'd156224;
    dina = {96'd0, 16'd4564, 16'd16904, 16'd57408, 16'd46661, 16'd65464, 16'd4159, 16'd20497, 16'd37927, 16'd19792, 16'd57270}; // indx = 4882
    #10;
    addra = 32'd156256;
    dina = {96'd0, 16'd24240, 16'd750, 16'd48079, 16'd63553, 16'd10011, 16'd53583, 16'd30410, 16'd15017, 16'd46324, 16'd2546}; // indx = 4883
    #10;
    addra = 32'd156288;
    dina = {96'd0, 16'd53072, 16'd58867, 16'd18299, 16'd5642, 16'd28028, 16'd28519, 16'd45522, 16'd34440, 16'd6379, 16'd26520}; // indx = 4884
    #10;
    addra = 32'd156320;
    dina = {96'd0, 16'd10650, 16'd38872, 16'd23701, 16'd25229, 16'd58832, 16'd50595, 16'd5506, 16'd49198, 16'd55323, 16'd7181}; // indx = 4885
    #10;
    addra = 32'd156352;
    dina = {96'd0, 16'd41173, 16'd5702, 16'd40265, 16'd43584, 16'd60354, 16'd20635, 16'd42338, 16'd30915, 16'd38355, 16'd65077}; // indx = 4886
    #10;
    addra = 32'd156384;
    dina = {96'd0, 16'd48288, 16'd12119, 16'd50254, 16'd6866, 16'd24449, 16'd28179, 16'd3837, 16'd64292, 16'd46316, 16'd59900}; // indx = 4887
    #10;
    addra = 32'd156416;
    dina = {96'd0, 16'd14885, 16'd58530, 16'd56498, 16'd16849, 16'd46817, 16'd16893, 16'd49929, 16'd27767, 16'd58729, 16'd50342}; // indx = 4888
    #10;
    addra = 32'd156448;
    dina = {96'd0, 16'd5889, 16'd45838, 16'd6514, 16'd51822, 16'd59786, 16'd27415, 16'd8311, 16'd42489, 16'd48580, 16'd4692}; // indx = 4889
    #10;
    addra = 32'd156480;
    dina = {96'd0, 16'd11755, 16'd52235, 16'd18960, 16'd64023, 16'd1950, 16'd62994, 16'd60543, 16'd38434, 16'd548, 16'd14651}; // indx = 4890
    #10;
    addra = 32'd156512;
    dina = {96'd0, 16'd42600, 16'd64408, 16'd54959, 16'd10999, 16'd8215, 16'd10882, 16'd36000, 16'd1508, 16'd8758, 16'd5383}; // indx = 4891
    #10;
    addra = 32'd156544;
    dina = {96'd0, 16'd63265, 16'd22878, 16'd61111, 16'd14548, 16'd19667, 16'd8749, 16'd64149, 16'd30879, 16'd9318, 16'd34136}; // indx = 4892
    #10;
    addra = 32'd156576;
    dina = {96'd0, 16'd45425, 16'd8365, 16'd30544, 16'd33115, 16'd998, 16'd13676, 16'd18061, 16'd32842, 16'd8926, 16'd61534}; // indx = 4893
    #10;
    addra = 32'd156608;
    dina = {96'd0, 16'd21989, 16'd54980, 16'd42135, 16'd62311, 16'd21527, 16'd4555, 16'd31741, 16'd41776, 16'd41441, 16'd46952}; // indx = 4894
    #10;
    addra = 32'd156640;
    dina = {96'd0, 16'd61571, 16'd34336, 16'd2421, 16'd48865, 16'd38505, 16'd13214, 16'd43767, 16'd18665, 16'd5744, 16'd17422}; // indx = 4895
    #10;
    addra = 32'd156672;
    dina = {96'd0, 16'd14203, 16'd34735, 16'd10845, 16'd41933, 16'd55389, 16'd14455, 16'd8515, 16'd21407, 16'd35985, 16'd46302}; // indx = 4896
    #10;
    addra = 32'd156704;
    dina = {96'd0, 16'd17328, 16'd52845, 16'd63475, 16'd48148, 16'd414, 16'd31075, 16'd13049, 16'd28214, 16'd40928, 16'd25563}; // indx = 4897
    #10;
    addra = 32'd156736;
    dina = {96'd0, 16'd1867, 16'd9428, 16'd52792, 16'd52440, 16'd35908, 16'd15939, 16'd37826, 16'd40548, 16'd2441, 16'd38617}; // indx = 4898
    #10;
    addra = 32'd156768;
    dina = {96'd0, 16'd44567, 16'd20921, 16'd44120, 16'd2511, 16'd60719, 16'd41798, 16'd25133, 16'd53685, 16'd5455, 16'd12679}; // indx = 4899
    #10;
    addra = 32'd156800;
    dina = {96'd0, 16'd13638, 16'd40588, 16'd61953, 16'd22464, 16'd17999, 16'd46780, 16'd5439, 16'd21585, 16'd33356, 16'd12956}; // indx = 4900
    #10;
    addra = 32'd156832;
    dina = {96'd0, 16'd36822, 16'd2809, 16'd42171, 16'd31371, 16'd279, 16'd27270, 16'd29053, 16'd12584, 16'd58904, 16'd63788}; // indx = 4901
    #10;
    addra = 32'd156864;
    dina = {96'd0, 16'd21913, 16'd64126, 16'd25715, 16'd32446, 16'd4208, 16'd50841, 16'd19272, 16'd36304, 16'd5699, 16'd45727}; // indx = 4902
    #10;
    addra = 32'd156896;
    dina = {96'd0, 16'd44253, 16'd54616, 16'd63791, 16'd18584, 16'd35783, 16'd26299, 16'd20293, 16'd57606, 16'd6881, 16'd26913}; // indx = 4903
    #10;
    addra = 32'd156928;
    dina = {96'd0, 16'd56240, 16'd37795, 16'd17646, 16'd31125, 16'd47749, 16'd25815, 16'd42026, 16'd43672, 16'd44085, 16'd34590}; // indx = 4904
    #10;
    addra = 32'd156960;
    dina = {96'd0, 16'd47014, 16'd20280, 16'd23443, 16'd48714, 16'd41874, 16'd1737, 16'd50178, 16'd26884, 16'd26036, 16'd20047}; // indx = 4905
    #10;
    addra = 32'd156992;
    dina = {96'd0, 16'd18523, 16'd55492, 16'd41637, 16'd13111, 16'd2755, 16'd60054, 16'd43614, 16'd19330, 16'd18980, 16'd53373}; // indx = 4906
    #10;
    addra = 32'd157024;
    dina = {96'd0, 16'd26073, 16'd54240, 16'd23796, 16'd44039, 16'd56810, 16'd28782, 16'd56532, 16'd7505, 16'd38663, 16'd31608}; // indx = 4907
    #10;
    addra = 32'd157056;
    dina = {96'd0, 16'd29461, 16'd27213, 16'd7694, 16'd47346, 16'd58652, 16'd60001, 16'd63960, 16'd43596, 16'd55828, 16'd64725}; // indx = 4908
    #10;
    addra = 32'd157088;
    dina = {96'd0, 16'd30948, 16'd24409, 16'd39233, 16'd48907, 16'd22878, 16'd25617, 16'd54549, 16'd7987, 16'd30861, 16'd40684}; // indx = 4909
    #10;
    addra = 32'd157120;
    dina = {96'd0, 16'd7761, 16'd20332, 16'd45625, 16'd2519, 16'd31634, 16'd51033, 16'd12449, 16'd34505, 16'd59488, 16'd63677}; // indx = 4910
    #10;
    addra = 32'd157152;
    dina = {96'd0, 16'd58772, 16'd19708, 16'd51195, 16'd29800, 16'd13856, 16'd23428, 16'd5933, 16'd9800, 16'd43413, 16'd62598}; // indx = 4911
    #10;
    addra = 32'd157184;
    dina = {96'd0, 16'd48625, 16'd49290, 16'd31133, 16'd10252, 16'd11405, 16'd17914, 16'd5519, 16'd54066, 16'd13451, 16'd11788}; // indx = 4912
    #10;
    addra = 32'd157216;
    dina = {96'd0, 16'd37380, 16'd64089, 16'd9302, 16'd31445, 16'd13113, 16'd57839, 16'd695, 16'd62244, 16'd64364, 16'd59137}; // indx = 4913
    #10;
    addra = 32'd157248;
    dina = {96'd0, 16'd36142, 16'd49499, 16'd30478, 16'd58176, 16'd50705, 16'd49601, 16'd21064, 16'd2253, 16'd36053, 16'd33540}; // indx = 4914
    #10;
    addra = 32'd157280;
    dina = {96'd0, 16'd40337, 16'd22257, 16'd22505, 16'd56374, 16'd1831, 16'd16279, 16'd53649, 16'd21756, 16'd1848, 16'd29228}; // indx = 4915
    #10;
    addra = 32'd157312;
    dina = {96'd0, 16'd50262, 16'd17960, 16'd30978, 16'd2623, 16'd19016, 16'd61823, 16'd42405, 16'd7068, 16'd6999, 16'd18869}; // indx = 4916
    #10;
    addra = 32'd157344;
    dina = {96'd0, 16'd10340, 16'd58546, 16'd6626, 16'd41902, 16'd4768, 16'd18788, 16'd53124, 16'd40127, 16'd22904, 16'd6574}; // indx = 4917
    #10;
    addra = 32'd157376;
    dina = {96'd0, 16'd34176, 16'd49376, 16'd41304, 16'd12055, 16'd8541, 16'd38612, 16'd29212, 16'd3677, 16'd23159, 16'd46196}; // indx = 4918
    #10;
    addra = 32'd157408;
    dina = {96'd0, 16'd49370, 16'd45124, 16'd14385, 16'd47840, 16'd28125, 16'd59186, 16'd31180, 16'd62164, 16'd39852, 16'd53517}; // indx = 4919
    #10;
    addra = 32'd157440;
    dina = {96'd0, 16'd2351, 16'd2280, 16'd14136, 16'd35194, 16'd45873, 16'd10723, 16'd43962, 16'd4791, 16'd59470, 16'd31589}; // indx = 4920
    #10;
    addra = 32'd157472;
    dina = {96'd0, 16'd28368, 16'd28429, 16'd30569, 16'd41155, 16'd15680, 16'd50531, 16'd14617, 16'd18007, 16'd24350, 16'd18187}; // indx = 4921
    #10;
    addra = 32'd157504;
    dina = {96'd0, 16'd44068, 16'd56261, 16'd606, 16'd23855, 16'd14194, 16'd25270, 16'd24005, 16'd50468, 16'd4368, 16'd41955}; // indx = 4922
    #10;
    addra = 32'd157536;
    dina = {96'd0, 16'd11512, 16'd7335, 16'd54679, 16'd5777, 16'd10340, 16'd26920, 16'd25855, 16'd10742, 16'd52277, 16'd56542}; // indx = 4923
    #10;
    addra = 32'd157568;
    dina = {96'd0, 16'd60657, 16'd24747, 16'd29236, 16'd42200, 16'd31425, 16'd62948, 16'd3670, 16'd51443, 16'd24512, 16'd13416}; // indx = 4924
    #10;
    addra = 32'd157600;
    dina = {96'd0, 16'd62086, 16'd33852, 16'd11839, 16'd63665, 16'd1225, 16'd44234, 16'd64892, 16'd11676, 16'd1968, 16'd16816}; // indx = 4925
    #10;
    addra = 32'd157632;
    dina = {96'd0, 16'd12100, 16'd26106, 16'd28402, 16'd39456, 16'd27612, 16'd41191, 16'd2375, 16'd6445, 16'd36259, 16'd41268}; // indx = 4926
    #10;
    addra = 32'd157664;
    dina = {96'd0, 16'd22795, 16'd44771, 16'd14435, 16'd4914, 16'd11352, 16'd63893, 16'd51439, 16'd35556, 16'd59626, 16'd48189}; // indx = 4927
    #10;
    addra = 32'd157696;
    dina = {96'd0, 16'd12179, 16'd6234, 16'd8050, 16'd15363, 16'd34631, 16'd38908, 16'd52001, 16'd55559, 16'd36252, 16'd11420}; // indx = 4928
    #10;
    addra = 32'd157728;
    dina = {96'd0, 16'd52199, 16'd61228, 16'd64358, 16'd51946, 16'd58043, 16'd15314, 16'd18723, 16'd3278, 16'd36627, 16'd53063}; // indx = 4929
    #10;
    addra = 32'd157760;
    dina = {96'd0, 16'd12943, 16'd4567, 16'd26399, 16'd60692, 16'd16046, 16'd45862, 16'd10390, 16'd48860, 16'd43774, 16'd33565}; // indx = 4930
    #10;
    addra = 32'd157792;
    dina = {96'd0, 16'd19411, 16'd16622, 16'd3109, 16'd50819, 16'd6289, 16'd37814, 16'd45457, 16'd52768, 16'd21805, 16'd48172}; // indx = 4931
    #10;
    addra = 32'd157824;
    dina = {96'd0, 16'd49136, 16'd7539, 16'd17133, 16'd42616, 16'd52049, 16'd32089, 16'd43613, 16'd7323, 16'd50648, 16'd53844}; // indx = 4932
    #10;
    addra = 32'd157856;
    dina = {96'd0, 16'd5200, 16'd17293, 16'd30356, 16'd16530, 16'd11841, 16'd64937, 16'd24547, 16'd29753, 16'd57488, 16'd28880}; // indx = 4933
    #10;
    addra = 32'd157888;
    dina = {96'd0, 16'd8138, 16'd60482, 16'd61646, 16'd62533, 16'd41183, 16'd58117, 16'd27266, 16'd39470, 16'd16767, 16'd54377}; // indx = 4934
    #10;
    addra = 32'd157920;
    dina = {96'd0, 16'd7619, 16'd36752, 16'd28510, 16'd819, 16'd40112, 16'd46550, 16'd1359, 16'd64742, 16'd22015, 16'd51310}; // indx = 4935
    #10;
    addra = 32'd157952;
    dina = {96'd0, 16'd33518, 16'd63253, 16'd17821, 16'd49475, 16'd31123, 16'd36862, 16'd53533, 16'd52041, 16'd21586, 16'd20291}; // indx = 4936
    #10;
    addra = 32'd157984;
    dina = {96'd0, 16'd59022, 16'd19505, 16'd36330, 16'd30502, 16'd16540, 16'd5647, 16'd4409, 16'd1865, 16'd34194, 16'd24519}; // indx = 4937
    #10;
    addra = 32'd158016;
    dina = {96'd0, 16'd58813, 16'd36538, 16'd57300, 16'd57645, 16'd33107, 16'd38521, 16'd65526, 16'd25556, 16'd3596, 16'd5795}; // indx = 4938
    #10;
    addra = 32'd158048;
    dina = {96'd0, 16'd37669, 16'd23595, 16'd55594, 16'd54074, 16'd63378, 16'd52559, 16'd40503, 16'd16673, 16'd9667, 16'd11377}; // indx = 4939
    #10;
    addra = 32'd158080;
    dina = {96'd0, 16'd50789, 16'd4222, 16'd48384, 16'd15203, 16'd34195, 16'd44759, 16'd42856, 16'd1608, 16'd58625, 16'd17836}; // indx = 4940
    #10;
    addra = 32'd158112;
    dina = {96'd0, 16'd59837, 16'd651, 16'd39287, 16'd5722, 16'd35119, 16'd52295, 16'd53711, 16'd46260, 16'd39376, 16'd53725}; // indx = 4941
    #10;
    addra = 32'd158144;
    dina = {96'd0, 16'd32241, 16'd26671, 16'd9636, 16'd16498, 16'd58592, 16'd31342, 16'd36554, 16'd9206, 16'd43705, 16'd49354}; // indx = 4942
    #10;
    addra = 32'd158176;
    dina = {96'd0, 16'd21575, 16'd63487, 16'd33557, 16'd50039, 16'd16330, 16'd37922, 16'd11346, 16'd29063, 16'd32438, 16'd37322}; // indx = 4943
    #10;
    addra = 32'd158208;
    dina = {96'd0, 16'd30833, 16'd3237, 16'd37931, 16'd8455, 16'd52394, 16'd58572, 16'd49074, 16'd63157, 16'd6011, 16'd49644}; // indx = 4944
    #10;
    addra = 32'd158240;
    dina = {96'd0, 16'd34874, 16'd25129, 16'd12509, 16'd42883, 16'd57820, 16'd45150, 16'd24820, 16'd29177, 16'd32430, 16'd62658}; // indx = 4945
    #10;
    addra = 32'd158272;
    dina = {96'd0, 16'd32604, 16'd31640, 16'd32625, 16'd14245, 16'd27052, 16'd40931, 16'd41872, 16'd62977, 16'd10236, 16'd64545}; // indx = 4946
    #10;
    addra = 32'd158304;
    dina = {96'd0, 16'd2772, 16'd34260, 16'd41657, 16'd33251, 16'd40509, 16'd16191, 16'd6091, 16'd42188, 16'd64156, 16'd15392}; // indx = 4947
    #10;
    addra = 32'd158336;
    dina = {96'd0, 16'd14699, 16'd23432, 16'd44774, 16'd4318, 16'd28350, 16'd44450, 16'd35633, 16'd14490, 16'd40284, 16'd36946}; // indx = 4948
    #10;
    addra = 32'd158368;
    dina = {96'd0, 16'd25506, 16'd25474, 16'd24532, 16'd25459, 16'd315, 16'd28654, 16'd2901, 16'd39297, 16'd36476, 16'd41871}; // indx = 4949
    #10;
    addra = 32'd158400;
    dina = {96'd0, 16'd63446, 16'd27927, 16'd11688, 16'd23191, 16'd64287, 16'd46795, 16'd20571, 16'd6915, 16'd6103, 16'd34168}; // indx = 4950
    #10;
    addra = 32'd158432;
    dina = {96'd0, 16'd13482, 16'd27027, 16'd2926, 16'd23601, 16'd17520, 16'd11570, 16'd64060, 16'd12139, 16'd55679, 16'd16019}; // indx = 4951
    #10;
    addra = 32'd158464;
    dina = {96'd0, 16'd30051, 16'd21396, 16'd61824, 16'd2201, 16'd33823, 16'd13961, 16'd59122, 16'd52589, 16'd30384, 16'd7011}; // indx = 4952
    #10;
    addra = 32'd158496;
    dina = {96'd0, 16'd19232, 16'd27776, 16'd18097, 16'd37937, 16'd14514, 16'd63229, 16'd18123, 16'd25777, 16'd16442, 16'd28906}; // indx = 4953
    #10;
    addra = 32'd158528;
    dina = {96'd0, 16'd30633, 16'd59364, 16'd12793, 16'd10033, 16'd14933, 16'd46292, 16'd52927, 16'd9062, 16'd35212, 16'd38043}; // indx = 4954
    #10;
    addra = 32'd158560;
    dina = {96'd0, 16'd33662, 16'd18519, 16'd8502, 16'd37612, 16'd20800, 16'd61456, 16'd11449, 16'd53135, 16'd45822, 16'd43592}; // indx = 4955
    #10;
    addra = 32'd158592;
    dina = {96'd0, 16'd18060, 16'd553, 16'd46492, 16'd58076, 16'd32608, 16'd45460, 16'd63908, 16'd40040, 16'd26570, 16'd41915}; // indx = 4956
    #10;
    addra = 32'd158624;
    dina = {96'd0, 16'd14452, 16'd23061, 16'd49172, 16'd2713, 16'd39529, 16'd13020, 16'd11375, 16'd25369, 16'd18051, 16'd41160}; // indx = 4957
    #10;
    addra = 32'd158656;
    dina = {96'd0, 16'd56730, 16'd55362, 16'd18672, 16'd46622, 16'd35921, 16'd46611, 16'd5175, 16'd4109, 16'd18288, 16'd30416}; // indx = 4958
    #10;
    addra = 32'd158688;
    dina = {96'd0, 16'd37110, 16'd37467, 16'd24305, 16'd4817, 16'd7066, 16'd55106, 16'd19607, 16'd42047, 16'd33445, 16'd48150}; // indx = 4959
    #10;
    addra = 32'd158720;
    dina = {96'd0, 16'd46296, 16'd61551, 16'd60082, 16'd64499, 16'd24122, 16'd47873, 16'd22097, 16'd30957, 16'd18428, 16'd54880}; // indx = 4960
    #10;
    addra = 32'd158752;
    dina = {96'd0, 16'd36402, 16'd454, 16'd11501, 16'd4247, 16'd44610, 16'd57972, 16'd49774, 16'd8578, 16'd6865, 16'd13398}; // indx = 4961
    #10;
    addra = 32'd158784;
    dina = {96'd0, 16'd18575, 16'd51763, 16'd62311, 16'd57465, 16'd13376, 16'd37602, 16'd14904, 16'd24003, 16'd6443, 16'd18839}; // indx = 4962
    #10;
    addra = 32'd158816;
    dina = {96'd0, 16'd50992, 16'd11729, 16'd56743, 16'd10390, 16'd16073, 16'd38450, 16'd13679, 16'd54039, 16'd55568, 16'd65498}; // indx = 4963
    #10;
    addra = 32'd158848;
    dina = {96'd0, 16'd37798, 16'd22630, 16'd54294, 16'd46258, 16'd34087, 16'd28617, 16'd50488, 16'd48293, 16'd47878, 16'd53784}; // indx = 4964
    #10;
    addra = 32'd158880;
    dina = {96'd0, 16'd32945, 16'd20155, 16'd31329, 16'd25307, 16'd35805, 16'd5243, 16'd7846, 16'd23168, 16'd64757, 16'd40787}; // indx = 4965
    #10;
    addra = 32'd158912;
    dina = {96'd0, 16'd62197, 16'd47815, 16'd10165, 16'd7911, 16'd17477, 16'd26096, 16'd27134, 16'd44330, 16'd6239, 16'd46460}; // indx = 4966
    #10;
    addra = 32'd158944;
    dina = {96'd0, 16'd24065, 16'd26849, 16'd95, 16'd34728, 16'd48663, 16'd56645, 16'd22125, 16'd13346, 16'd6437, 16'd60051}; // indx = 4967
    #10;
    addra = 32'd158976;
    dina = {96'd0, 16'd55691, 16'd24182, 16'd20111, 16'd56447, 16'd52814, 16'd33434, 16'd18471, 16'd48111, 16'd52157, 16'd49853}; // indx = 4968
    #10;
    addra = 32'd159008;
    dina = {96'd0, 16'd31893, 16'd16788, 16'd40584, 16'd17727, 16'd22538, 16'd31540, 16'd28343, 16'd26005, 16'd38627, 16'd21051}; // indx = 4969
    #10;
    addra = 32'd159040;
    dina = {96'd0, 16'd49679, 16'd50800, 16'd25947, 16'd29398, 16'd65322, 16'd23283, 16'd64698, 16'd35389, 16'd19955, 16'd62775}; // indx = 4970
    #10;
    addra = 32'd159072;
    dina = {96'd0, 16'd54124, 16'd35252, 16'd6323, 16'd60481, 16'd37114, 16'd52102, 16'd9977, 16'd47555, 16'd511, 16'd31285}; // indx = 4971
    #10;
    addra = 32'd159104;
    dina = {96'd0, 16'd22792, 16'd38297, 16'd33349, 16'd54490, 16'd36666, 16'd41659, 16'd2322, 16'd51304, 16'd19221, 16'd53102}; // indx = 4972
    #10;
    addra = 32'd159136;
    dina = {96'd0, 16'd48864, 16'd39220, 16'd16768, 16'd19044, 16'd9618, 16'd18402, 16'd52296, 16'd19475, 16'd51088, 16'd53085}; // indx = 4973
    #10;
    addra = 32'd159168;
    dina = {96'd0, 16'd33287, 16'd47058, 16'd41357, 16'd3863, 16'd23747, 16'd15241, 16'd45450, 16'd57446, 16'd49305, 16'd33751}; // indx = 4974
    #10;
    addra = 32'd159200;
    dina = {96'd0, 16'd59550, 16'd6526, 16'd2176, 16'd7810, 16'd11557, 16'd48906, 16'd64505, 16'd44588, 16'd56252, 16'd20269}; // indx = 4975
    #10;
    addra = 32'd159232;
    dina = {96'd0, 16'd53135, 16'd13453, 16'd34424, 16'd44547, 16'd58480, 16'd36979, 16'd44636, 16'd34019, 16'd15538, 16'd29642}; // indx = 4976
    #10;
    addra = 32'd159264;
    dina = {96'd0, 16'd36658, 16'd60140, 16'd20011, 16'd5165, 16'd47242, 16'd29690, 16'd16837, 16'd21863, 16'd740, 16'd8920}; // indx = 4977
    #10;
    addra = 32'd159296;
    dina = {96'd0, 16'd61420, 16'd44382, 16'd65203, 16'd33335, 16'd40706, 16'd13421, 16'd29642, 16'd13527, 16'd41256, 16'd39811}; // indx = 4978
    #10;
    addra = 32'd159328;
    dina = {96'd0, 16'd63672, 16'd30694, 16'd54373, 16'd42280, 16'd32297, 16'd56882, 16'd49262, 16'd33476, 16'd31450, 16'd49504}; // indx = 4979
    #10;
    addra = 32'd159360;
    dina = {96'd0, 16'd2279, 16'd1973, 16'd34373, 16'd57322, 16'd10090, 16'd27082, 16'd28030, 16'd36096, 16'd62658, 16'd19291}; // indx = 4980
    #10;
    addra = 32'd159392;
    dina = {96'd0, 16'd55638, 16'd44101, 16'd38951, 16'd36544, 16'd33854, 16'd42726, 16'd9180, 16'd41890, 16'd19467, 16'd10486}; // indx = 4981
    #10;
    addra = 32'd159424;
    dina = {96'd0, 16'd65258, 16'd47537, 16'd355, 16'd20885, 16'd18690, 16'd46542, 16'd2448, 16'd40727, 16'd5942, 16'd57522}; // indx = 4982
    #10;
    addra = 32'd159456;
    dina = {96'd0, 16'd37969, 16'd53571, 16'd45995, 16'd24117, 16'd34669, 16'd46214, 16'd7790, 16'd24293, 16'd60225, 16'd34377}; // indx = 4983
    #10;
    addra = 32'd159488;
    dina = {96'd0, 16'd33804, 16'd34659, 16'd1993, 16'd39742, 16'd8732, 16'd61140, 16'd47686, 16'd25007, 16'd17126, 16'd26444}; // indx = 4984
    #10;
    addra = 32'd159520;
    dina = {96'd0, 16'd19215, 16'd32608, 16'd5485, 16'd9190, 16'd55063, 16'd48807, 16'd11559, 16'd4685, 16'd31023, 16'd57614}; // indx = 4985
    #10;
    addra = 32'd159552;
    dina = {96'd0, 16'd44953, 16'd63931, 16'd14848, 16'd1242, 16'd27629, 16'd61190, 16'd3585, 16'd40161, 16'd25377, 16'd37328}; // indx = 4986
    #10;
    addra = 32'd159584;
    dina = {96'd0, 16'd50945, 16'd37047, 16'd7298, 16'd55551, 16'd59648, 16'd8089, 16'd59490, 16'd4078, 16'd25132, 16'd21690}; // indx = 4987
    #10;
    addra = 32'd159616;
    dina = {96'd0, 16'd23697, 16'd38191, 16'd54291, 16'd38854, 16'd36737, 16'd41248, 16'd24248, 16'd11617, 16'd31350, 16'd55434}; // indx = 4988
    #10;
    addra = 32'd159648;
    dina = {96'd0, 16'd64062, 16'd24128, 16'd31600, 16'd45790, 16'd11065, 16'd272, 16'd46977, 16'd34219, 16'd5922, 16'd18852}; // indx = 4989
    #10;
    addra = 32'd159680;
    dina = {96'd0, 16'd34609, 16'd3573, 16'd58002, 16'd703, 16'd53589, 16'd49787, 16'd23500, 16'd29711, 16'd8228, 16'd40862}; // indx = 4990
    #10;
    addra = 32'd159712;
    dina = {96'd0, 16'd17404, 16'd37284, 16'd36711, 16'd18778, 16'd35026, 16'd18397, 16'd47002, 16'd59808, 16'd52883, 16'd47268}; // indx = 4991
    #10;
    addra = 32'd159744;
    dina = {96'd0, 16'd55267, 16'd64029, 16'd22541, 16'd29251, 16'd15721, 16'd52913, 16'd43139, 16'd39470, 16'd34233, 16'd62883}; // indx = 4992
    #10;
    addra = 32'd159776;
    dina = {96'd0, 16'd36695, 16'd28370, 16'd9332, 16'd5734, 16'd45044, 16'd15643, 16'd18148, 16'd29366, 16'd22517, 16'd64787}; // indx = 4993
    #10;
    addra = 32'd159808;
    dina = {96'd0, 16'd14705, 16'd37097, 16'd59360, 16'd39883, 16'd24042, 16'd20919, 16'd45758, 16'd26710, 16'd13837, 16'd6222}; // indx = 4994
    #10;
    addra = 32'd159840;
    dina = {96'd0, 16'd51667, 16'd58193, 16'd28476, 16'd49051, 16'd19540, 16'd62804, 16'd555, 16'd7124, 16'd52795, 16'd63480}; // indx = 4995
    #10;
    addra = 32'd159872;
    dina = {96'd0, 16'd38135, 16'd10931, 16'd56720, 16'd40826, 16'd858, 16'd37767, 16'd1764, 16'd1554, 16'd42314, 16'd11415}; // indx = 4996
    #10;
    addra = 32'd159904;
    dina = {96'd0, 16'd9055, 16'd27621, 16'd8841, 16'd17651, 16'd51013, 16'd1789, 16'd57811, 16'd29337, 16'd21972, 16'd61065}; // indx = 4997
    #10;
    addra = 32'd159936;
    dina = {96'd0, 16'd27067, 16'd14401, 16'd14594, 16'd23943, 16'd11966, 16'd52673, 16'd48543, 16'd17309, 16'd63676, 16'd52075}; // indx = 4998
    #10;
    addra = 32'd159968;
    dina = {96'd0, 16'd10186, 16'd60665, 16'd28365, 16'd26769, 16'd17526, 16'd59154, 16'd42399, 16'd60832, 16'd19409, 16'd42083}; // indx = 4999
    #10;
    addra = 32'd160000;
    dina = {96'd0, 16'd4092, 16'd41914, 16'd31876, 16'd19603, 16'd2790, 16'd40883, 16'd22323, 16'd54439, 16'd33847, 16'd62504}; // indx = 5000
    #10;
    addra = 32'd160032;
    dina = {96'd0, 16'd14963, 16'd4522, 16'd26615, 16'd16501, 16'd63358, 16'd45843, 16'd4057, 16'd6118, 16'd25632, 16'd3652}; // indx = 5001
    #10;
    addra = 32'd160064;
    dina = {96'd0, 16'd23958, 16'd48979, 16'd63695, 16'd33887, 16'd27811, 16'd54048, 16'd47240, 16'd57236, 16'd37421, 16'd30912}; // indx = 5002
    #10;
    addra = 32'd160096;
    dina = {96'd0, 16'd31926, 16'd11750, 16'd7932, 16'd24536, 16'd43799, 16'd25694, 16'd56392, 16'd43240, 16'd40696, 16'd15181}; // indx = 5003
    #10;
    addra = 32'd160128;
    dina = {96'd0, 16'd27985, 16'd51209, 16'd3316, 16'd62732, 16'd959, 16'd32512, 16'd26284, 16'd9265, 16'd47719, 16'd29995}; // indx = 5004
    #10;
    addra = 32'd160160;
    dina = {96'd0, 16'd25389, 16'd60225, 16'd60070, 16'd55303, 16'd50871, 16'd21222, 16'd43784, 16'd53523, 16'd29222, 16'd59161}; // indx = 5005
    #10;
    addra = 32'd160192;
    dina = {96'd0, 16'd41763, 16'd9105, 16'd11788, 16'd2319, 16'd46619, 16'd36938, 16'd64988, 16'd22522, 16'd7995, 16'd47184}; // indx = 5006
    #10;
    addra = 32'd160224;
    dina = {96'd0, 16'd47412, 16'd51838, 16'd61000, 16'd7341, 16'd46047, 16'd31287, 16'd59599, 16'd58887, 16'd36023, 16'd13092}; // indx = 5007
    #10;
    addra = 32'd160256;
    dina = {96'd0, 16'd50152, 16'd25882, 16'd46114, 16'd20818, 16'd46325, 16'd7333, 16'd9028, 16'd14331, 16'd20305, 16'd31054}; // indx = 5008
    #10;
    addra = 32'd160288;
    dina = {96'd0, 16'd11924, 16'd37231, 16'd53403, 16'd4704, 16'd6287, 16'd15969, 16'd51, 16'd29944, 16'd41916, 16'd220}; // indx = 5009
    #10;
    addra = 32'd160320;
    dina = {96'd0, 16'd39607, 16'd40608, 16'd42932, 16'd1437, 16'd37609, 16'd5312, 16'd59501, 16'd12766, 16'd4763, 16'd20314}; // indx = 5010
    #10;
    addra = 32'd160352;
    dina = {96'd0, 16'd7446, 16'd8936, 16'd37278, 16'd17263, 16'd989, 16'd16306, 16'd30821, 16'd26079, 16'd21973, 16'd65138}; // indx = 5011
    #10;
    addra = 32'd160384;
    dina = {96'd0, 16'd30097, 16'd38917, 16'd10346, 16'd47045, 16'd24411, 16'd49003, 16'd22008, 16'd6713, 16'd51653, 16'd14724}; // indx = 5012
    #10;
    addra = 32'd160416;
    dina = {96'd0, 16'd19973, 16'd16841, 16'd32528, 16'd18228, 16'd8506, 16'd48513, 16'd62044, 16'd54727, 16'd36902, 16'd41136}; // indx = 5013
    #10;
    addra = 32'd160448;
    dina = {96'd0, 16'd20953, 16'd58372, 16'd31518, 16'd39409, 16'd8078, 16'd38858, 16'd41410, 16'd60253, 16'd63900, 16'd19987}; // indx = 5014
    #10;
    addra = 32'd160480;
    dina = {96'd0, 16'd48654, 16'd48599, 16'd26206, 16'd47589, 16'd33407, 16'd15349, 16'd59752, 16'd54001, 16'd60815, 16'd17673}; // indx = 5015
    #10;
    addra = 32'd160512;
    dina = {96'd0, 16'd35954, 16'd46635, 16'd37205, 16'd7930, 16'd20478, 16'd34546, 16'd10069, 16'd30965, 16'd43012, 16'd32443}; // indx = 5016
    #10;
    addra = 32'd160544;
    dina = {96'd0, 16'd52507, 16'd46202, 16'd31827, 16'd52687, 16'd46315, 16'd49187, 16'd25142, 16'd16015, 16'd29015, 16'd46390}; // indx = 5017
    #10;
    addra = 32'd160576;
    dina = {96'd0, 16'd48885, 16'd17761, 16'd53259, 16'd13998, 16'd27513, 16'd29458, 16'd20381, 16'd38139, 16'd44336, 16'd39021}; // indx = 5018
    #10;
    addra = 32'd160608;
    dina = {96'd0, 16'd17220, 16'd50411, 16'd28720, 16'd6600, 16'd54699, 16'd47888, 16'd38919, 16'd61897, 16'd42601, 16'd26526}; // indx = 5019
    #10;
    addra = 32'd160640;
    dina = {96'd0, 16'd11221, 16'd30666, 16'd2389, 16'd2375, 16'd2327, 16'd18019, 16'd26067, 16'd59913, 16'd1644, 16'd18933}; // indx = 5020
    #10;
    addra = 32'd160672;
    dina = {96'd0, 16'd21012, 16'd55147, 16'd61342, 16'd49917, 16'd27328, 16'd8597, 16'd39093, 16'd43900, 16'd17570, 16'd32275}; // indx = 5021
    #10;
    addra = 32'd160704;
    dina = {96'd0, 16'd14215, 16'd23106, 16'd58935, 16'd49504, 16'd31841, 16'd32914, 16'd56582, 16'd58138, 16'd29917, 16'd32749}; // indx = 5022
    #10;
    addra = 32'd160736;
    dina = {96'd0, 16'd22279, 16'd48465, 16'd54595, 16'd21795, 16'd43570, 16'd2063, 16'd29016, 16'd53539, 16'd26025, 16'd434}; // indx = 5023
    #10;
    addra = 32'd160768;
    dina = {96'd0, 16'd40894, 16'd42236, 16'd44368, 16'd46252, 16'd22898, 16'd35628, 16'd49445, 16'd36635, 16'd14235, 16'd57517}; // indx = 5024
    #10;
    addra = 32'd160800;
    dina = {96'd0, 16'd7026, 16'd39541, 16'd31643, 16'd58770, 16'd34376, 16'd5661, 16'd35924, 16'd12681, 16'd43939, 16'd49583}; // indx = 5025
    #10;
    addra = 32'd160832;
    dina = {96'd0, 16'd42594, 16'd8035, 16'd1330, 16'd44302, 16'd36916, 16'd9688, 16'd3567, 16'd12337, 16'd15589, 16'd48615}; // indx = 5026
    #10;
    addra = 32'd160864;
    dina = {96'd0, 16'd42742, 16'd41536, 16'd42770, 16'd59303, 16'd46595, 16'd21768, 16'd5556, 16'd61153, 16'd40222, 16'd39732}; // indx = 5027
    #10;
    addra = 32'd160896;
    dina = {96'd0, 16'd10169, 16'd34439, 16'd56994, 16'd61244, 16'd1888, 16'd65088, 16'd20119, 16'd52830, 16'd43679, 16'd39909}; // indx = 5028
    #10;
    addra = 32'd160928;
    dina = {96'd0, 16'd10874, 16'd996, 16'd38801, 16'd13269, 16'd60570, 16'd22684, 16'd62329, 16'd56065, 16'd22764, 16'd16088}; // indx = 5029
    #10;
    addra = 32'd160960;
    dina = {96'd0, 16'd48716, 16'd19227, 16'd50836, 16'd27298, 16'd54355, 16'd34740, 16'd8845, 16'd18510, 16'd26882, 16'd23391}; // indx = 5030
    #10;
    addra = 32'd160992;
    dina = {96'd0, 16'd1257, 16'd33488, 16'd27647, 16'd15818, 16'd47328, 16'd1550, 16'd11420, 16'd53616, 16'd53524, 16'd4978}; // indx = 5031
    #10;
    addra = 32'd161024;
    dina = {96'd0, 16'd15327, 16'd3395, 16'd18635, 16'd46034, 16'd5841, 16'd424, 16'd39402, 16'd46822, 16'd43150, 16'd61777}; // indx = 5032
    #10;
    addra = 32'd161056;
    dina = {96'd0, 16'd34726, 16'd35674, 16'd38108, 16'd2183, 16'd32305, 16'd5045, 16'd21735, 16'd51810, 16'd51281, 16'd24275}; // indx = 5033
    #10;
    addra = 32'd161088;
    dina = {96'd0, 16'd16459, 16'd61244, 16'd62014, 16'd62361, 16'd8016, 16'd18737, 16'd29136, 16'd65219, 16'd27903, 16'd44705}; // indx = 5034
    #10;
    addra = 32'd161120;
    dina = {96'd0, 16'd39416, 16'd14029, 16'd11049, 16'd9851, 16'd32420, 16'd43347, 16'd50285, 16'd28178, 16'd22629, 16'd14160}; // indx = 5035
    #10;
    addra = 32'd161152;
    dina = {96'd0, 16'd44467, 16'd32240, 16'd58089, 16'd13387, 16'd36387, 16'd53976, 16'd38411, 16'd24592, 16'd29187, 16'd34346}; // indx = 5036
    #10;
    addra = 32'd161184;
    dina = {96'd0, 16'd26302, 16'd3782, 16'd36440, 16'd10412, 16'd51137, 16'd59788, 16'd51131, 16'd55222, 16'd11796, 16'd64142}; // indx = 5037
    #10;
    addra = 32'd161216;
    dina = {96'd0, 16'd38735, 16'd31269, 16'd8940, 16'd13648, 16'd38351, 16'd12808, 16'd16223, 16'd39551, 16'd44750, 16'd2099}; // indx = 5038
    #10;
    addra = 32'd161248;
    dina = {96'd0, 16'd28091, 16'd11060, 16'd33334, 16'd32015, 16'd31491, 16'd27535, 16'd9281, 16'd2707, 16'd3044, 16'd31905}; // indx = 5039
    #10;
    addra = 32'd161280;
    dina = {96'd0, 16'd17949, 16'd55546, 16'd38654, 16'd14431, 16'd45120, 16'd64186, 16'd24397, 16'd57436, 16'd56100, 16'd12633}; // indx = 5040
    #10;
    addra = 32'd161312;
    dina = {96'd0, 16'd9603, 16'd64356, 16'd21758, 16'd62896, 16'd21536, 16'd56020, 16'd43890, 16'd36352, 16'd57730, 16'd3981}; // indx = 5041
    #10;
    addra = 32'd161344;
    dina = {96'd0, 16'd34678, 16'd20103, 16'd52817, 16'd4130, 16'd59751, 16'd52026, 16'd47295, 16'd8280, 16'd31461, 16'd14718}; // indx = 5042
    #10;
    addra = 32'd161376;
    dina = {96'd0, 16'd63269, 16'd15194, 16'd29806, 16'd20239, 16'd63216, 16'd48408, 16'd37765, 16'd24878, 16'd42415, 16'd7222}; // indx = 5043
    #10;
    addra = 32'd161408;
    dina = {96'd0, 16'd24413, 16'd8592, 16'd42541, 16'd60176, 16'd59481, 16'd49020, 16'd7237, 16'd52727, 16'd38, 16'd30920}; // indx = 5044
    #10;
    addra = 32'd161440;
    dina = {96'd0, 16'd29649, 16'd46325, 16'd44741, 16'd10395, 16'd49524, 16'd13473, 16'd18507, 16'd1625, 16'd7783, 16'd29831}; // indx = 5045
    #10;
    addra = 32'd161472;
    dina = {96'd0, 16'd37274, 16'd19425, 16'd23705, 16'd49695, 16'd13747, 16'd62889, 16'd35560, 16'd16268, 16'd33605, 16'd4055}; // indx = 5046
    #10;
    addra = 32'd161504;
    dina = {96'd0, 16'd56719, 16'd53379, 16'd24290, 16'd64229, 16'd37811, 16'd35459, 16'd19391, 16'd6395, 16'd23389, 16'd24368}; // indx = 5047
    #10;
    addra = 32'd161536;
    dina = {96'd0, 16'd41891, 16'd43052, 16'd19594, 16'd27235, 16'd28653, 16'd26444, 16'd31265, 16'd49136, 16'd28559, 16'd58217}; // indx = 5048
    #10;
    addra = 32'd161568;
    dina = {96'd0, 16'd3585, 16'd14158, 16'd36444, 16'd44904, 16'd8662, 16'd10680, 16'd45502, 16'd60992, 16'd35712, 16'd1022}; // indx = 5049
    #10;
    addra = 32'd161600;
    dina = {96'd0, 16'd21006, 16'd56266, 16'd54179, 16'd11835, 16'd13459, 16'd65522, 16'd15259, 16'd64990, 16'd25283, 16'd23820}; // indx = 5050
    #10;
    addra = 32'd161632;
    dina = {96'd0, 16'd33548, 16'd38445, 16'd24613, 16'd42557, 16'd60697, 16'd13833, 16'd8947, 16'd28359, 16'd27976, 16'd43951}; // indx = 5051
    #10;
    addra = 32'd161664;
    dina = {96'd0, 16'd20601, 16'd7427, 16'd16545, 16'd61193, 16'd34272, 16'd14978, 16'd61342, 16'd38002, 16'd19059, 16'd10343}; // indx = 5052
    #10;
    addra = 32'd161696;
    dina = {96'd0, 16'd151, 16'd28744, 16'd20779, 16'd53262, 16'd45814, 16'd63289, 16'd23709, 16'd57629, 16'd8740, 16'd13926}; // indx = 5053
    #10;
    addra = 32'd161728;
    dina = {96'd0, 16'd50703, 16'd18848, 16'd45073, 16'd4400, 16'd22572, 16'd19706, 16'd27197, 16'd22615, 16'd45470, 16'd5418}; // indx = 5054
    #10;
    addra = 32'd161760;
    dina = {96'd0, 16'd15896, 16'd27795, 16'd52176, 16'd65094, 16'd50746, 16'd58500, 16'd3556, 16'd56517, 16'd17698, 16'd33160}; // indx = 5055
    #10;
    addra = 32'd161792;
    dina = {96'd0, 16'd27565, 16'd34570, 16'd12074, 16'd25858, 16'd26440, 16'd59560, 16'd12836, 16'd47881, 16'd11624, 16'd47404}; // indx = 5056
    #10;
    addra = 32'd161824;
    dina = {96'd0, 16'd9789, 16'd61364, 16'd12754, 16'd65246, 16'd26365, 16'd23708, 16'd457, 16'd41951, 16'd45309, 16'd35659}; // indx = 5057
    #10;
    addra = 32'd161856;
    dina = {96'd0, 16'd1340, 16'd58379, 16'd20158, 16'd49954, 16'd41869, 16'd30810, 16'd33169, 16'd48067, 16'd57910, 16'd33267}; // indx = 5058
    #10;
    addra = 32'd161888;
    dina = {96'd0, 16'd5337, 16'd1174, 16'd62696, 16'd44787, 16'd7998, 16'd64403, 16'd44334, 16'd60203, 16'd18743, 16'd45365}; // indx = 5059
    #10;
    addra = 32'd161920;
    dina = {96'd0, 16'd9826, 16'd13480, 16'd41673, 16'd55474, 16'd37815, 16'd14568, 16'd27566, 16'd57250, 16'd7489, 16'd40486}; // indx = 5060
    #10;
    addra = 32'd161952;
    dina = {96'd0, 16'd55733, 16'd6592, 16'd37762, 16'd38825, 16'd53958, 16'd41886, 16'd50559, 16'd15055, 16'd51461, 16'd37530}; // indx = 5061
    #10;
    addra = 32'd161984;
    dina = {96'd0, 16'd35227, 16'd32720, 16'd44993, 16'd57446, 16'd11183, 16'd10749, 16'd34700, 16'd13658, 16'd22193, 16'd43636}; // indx = 5062
    #10;
    addra = 32'd162016;
    dina = {96'd0, 16'd14739, 16'd53648, 16'd48919, 16'd22411, 16'd52620, 16'd55230, 16'd19300, 16'd58904, 16'd61736, 16'd57461}; // indx = 5063
    #10;
    addra = 32'd162048;
    dina = {96'd0, 16'd24340, 16'd22433, 16'd12890, 16'd31280, 16'd54804, 16'd15757, 16'd35850, 16'd42312, 16'd64481, 16'd35463}; // indx = 5064
    #10;
    addra = 32'd162080;
    dina = {96'd0, 16'd50582, 16'd20104, 16'd43390, 16'd22824, 16'd36487, 16'd14986, 16'd30663, 16'd44962, 16'd21721, 16'd45891}; // indx = 5065
    #10;
    addra = 32'd162112;
    dina = {96'd0, 16'd25458, 16'd18270, 16'd42139, 16'd32230, 16'd8107, 16'd48447, 16'd1794, 16'd4413, 16'd13211, 16'd46374}; // indx = 5066
    #10;
    addra = 32'd162144;
    dina = {96'd0, 16'd64435, 16'd55000, 16'd11248, 16'd38199, 16'd50599, 16'd20589, 16'd63698, 16'd42588, 16'd27001, 16'd45918}; // indx = 5067
    #10;
    addra = 32'd162176;
    dina = {96'd0, 16'd13967, 16'd60994, 16'd38711, 16'd621, 16'd43022, 16'd27763, 16'd32126, 16'd52960, 16'd19957, 16'd24475}; // indx = 5068
    #10;
    addra = 32'd162208;
    dina = {96'd0, 16'd10091, 16'd3671, 16'd44018, 16'd54699, 16'd19946, 16'd40967, 16'd18280, 16'd9631, 16'd14206, 16'd43497}; // indx = 5069
    #10;
    addra = 32'd162240;
    dina = {96'd0, 16'd61559, 16'd36561, 16'd62941, 16'd42864, 16'd38929, 16'd61898, 16'd4136, 16'd60927, 16'd41313, 16'd36404}; // indx = 5070
    #10;
    addra = 32'd162272;
    dina = {96'd0, 16'd44852, 16'd55516, 16'd64830, 16'd18019, 16'd50375, 16'd15754, 16'd49905, 16'd62550, 16'd1397, 16'd23052}; // indx = 5071
    #10;
    addra = 32'd162304;
    dina = {96'd0, 16'd59715, 16'd34449, 16'd31474, 16'd18501, 16'd8897, 16'd53752, 16'd51384, 16'd61146, 16'd26293, 16'd3227}; // indx = 5072
    #10;
    addra = 32'd162336;
    dina = {96'd0, 16'd30129, 16'd852, 16'd20108, 16'd31288, 16'd52664, 16'd26642, 16'd38198, 16'd38637, 16'd34978, 16'd52171}; // indx = 5073
    #10;
    addra = 32'd162368;
    dina = {96'd0, 16'd38928, 16'd46843, 16'd17290, 16'd5921, 16'd58457, 16'd39073, 16'd14525, 16'd48229, 16'd18001, 16'd44852}; // indx = 5074
    #10;
    addra = 32'd162400;
    dina = {96'd0, 16'd11330, 16'd21612, 16'd4502, 16'd13918, 16'd52007, 16'd19114, 16'd56696, 16'd17891, 16'd50946, 16'd22924}; // indx = 5075
    #10;
    addra = 32'd162432;
    dina = {96'd0, 16'd25102, 16'd28849, 16'd42890, 16'd14065, 16'd31368, 16'd15553, 16'd30294, 16'd43369, 16'd15578, 16'd19494}; // indx = 5076
    #10;
    addra = 32'd162464;
    dina = {96'd0, 16'd45293, 16'd8797, 16'd19336, 16'd30953, 16'd63253, 16'd30666, 16'd62798, 16'd65263, 16'd6364, 16'd49806}; // indx = 5077
    #10;
    addra = 32'd162496;
    dina = {96'd0, 16'd47476, 16'd11044, 16'd35635, 16'd16180, 16'd60586, 16'd12009, 16'd48664, 16'd42471, 16'd61766, 16'd58348}; // indx = 5078
    #10;
    addra = 32'd162528;
    dina = {96'd0, 16'd29067, 16'd64441, 16'd60454, 16'd12266, 16'd14502, 16'd1567, 16'd19697, 16'd30621, 16'd2848, 16'd52967}; // indx = 5079
    #10;
    addra = 32'd162560;
    dina = {96'd0, 16'd30636, 16'd43672, 16'd6028, 16'd50039, 16'd61723, 16'd24725, 16'd15179, 16'd20424, 16'd63937, 16'd49959}; // indx = 5080
    #10;
    addra = 32'd162592;
    dina = {96'd0, 16'd10068, 16'd51205, 16'd7876, 16'd41645, 16'd48224, 16'd22627, 16'd1043, 16'd51945, 16'd50824, 16'd45426}; // indx = 5081
    #10;
    addra = 32'd162624;
    dina = {96'd0, 16'd52321, 16'd36171, 16'd33953, 16'd8913, 16'd50339, 16'd45208, 16'd64508, 16'd33203, 16'd29268, 16'd39602}; // indx = 5082
    #10;
    addra = 32'd162656;
    dina = {96'd0, 16'd58287, 16'd52023, 16'd23319, 16'd31349, 16'd58109, 16'd17199, 16'd38017, 16'd58843, 16'd39322, 16'd15775}; // indx = 5083
    #10;
    addra = 32'd162688;
    dina = {96'd0, 16'd13066, 16'd18231, 16'd57821, 16'd50767, 16'd45743, 16'd3864, 16'd4128, 16'd54751, 16'd61635, 16'd10405}; // indx = 5084
    #10;
    addra = 32'd162720;
    dina = {96'd0, 16'd29601, 16'd62117, 16'd53411, 16'd26267, 16'd6958, 16'd6134, 16'd24023, 16'd61503, 16'd22161, 16'd44037}; // indx = 5085
    #10;
    addra = 32'd162752;
    dina = {96'd0, 16'd18226, 16'd50729, 16'd50192, 16'd3614, 16'd61950, 16'd19055, 16'd16523, 16'd62241, 16'd13260, 16'd29639}; // indx = 5086
    #10;
    addra = 32'd162784;
    dina = {96'd0, 16'd36108, 16'd40999, 16'd36221, 16'd723, 16'd41309, 16'd40691, 16'd53735, 16'd5342, 16'd35639, 16'd51675}; // indx = 5087
    #10;
    addra = 32'd162816;
    dina = {96'd0, 16'd55957, 16'd4822, 16'd49031, 16'd56781, 16'd12559, 16'd38233, 16'd29078, 16'd37173, 16'd54711, 16'd47069}; // indx = 5088
    #10;
    addra = 32'd162848;
    dina = {96'd0, 16'd56712, 16'd22745, 16'd32077, 16'd54022, 16'd29718, 16'd41425, 16'd54297, 16'd30655, 16'd49913, 16'd26510}; // indx = 5089
    #10;
    addra = 32'd162880;
    dina = {96'd0, 16'd3563, 16'd2476, 16'd41855, 16'd5614, 16'd62728, 16'd24794, 16'd41742, 16'd55453, 16'd57186, 16'd51130}; // indx = 5090
    #10;
    addra = 32'd162912;
    dina = {96'd0, 16'd19263, 16'd48447, 16'd22733, 16'd3644, 16'd12128, 16'd57288, 16'd62354, 16'd4834, 16'd21469, 16'd25196}; // indx = 5091
    #10;
    addra = 32'd162944;
    dina = {96'd0, 16'd56593, 16'd48285, 16'd39509, 16'd16648, 16'd45202, 16'd4712, 16'd58316, 16'd50236, 16'd13313, 16'd15325}; // indx = 5092
    #10;
    addra = 32'd162976;
    dina = {96'd0, 16'd29756, 16'd28359, 16'd18447, 16'd38822, 16'd2964, 16'd60251, 16'd19315, 16'd12859, 16'd23544, 16'd12432}; // indx = 5093
    #10;
    addra = 32'd163008;
    dina = {96'd0, 16'd20810, 16'd48259, 16'd54372, 16'd18083, 16'd8613, 16'd7935, 16'd12649, 16'd43832, 16'd48906, 16'd57851}; // indx = 5094
    #10;
    addra = 32'd163040;
    dina = {96'd0, 16'd52999, 16'd59584, 16'd57715, 16'd26336, 16'd45976, 16'd3706, 16'd50811, 16'd6449, 16'd64403, 16'd15418}; // indx = 5095
    #10;
    addra = 32'd163072;
    dina = {96'd0, 16'd43132, 16'd19963, 16'd55309, 16'd49568, 16'd21650, 16'd15822, 16'd47315, 16'd13776, 16'd24501, 16'd6391}; // indx = 5096
    #10;
    addra = 32'd163104;
    dina = {96'd0, 16'd17442, 16'd37088, 16'd53567, 16'd8423, 16'd42626, 16'd24257, 16'd23425, 16'd40924, 16'd4240, 16'd24704}; // indx = 5097
    #10;
    addra = 32'd163136;
    dina = {96'd0, 16'd40355, 16'd11267, 16'd28492, 16'd23608, 16'd27403, 16'd54623, 16'd28452, 16'd17918, 16'd62667, 16'd63528}; // indx = 5098
    #10;
    addra = 32'd163168;
    dina = {96'd0, 16'd18562, 16'd41449, 16'd61754, 16'd54214, 16'd25920, 16'd32203, 16'd51500, 16'd17542, 16'd50710, 16'd54104}; // indx = 5099
    #10;
    addra = 32'd163200;
    dina = {96'd0, 16'd39657, 16'd15504, 16'd38813, 16'd5033, 16'd39403, 16'd43768, 16'd65009, 16'd60491, 16'd62224, 16'd58432}; // indx = 5100
    #10;
    addra = 32'd163232;
    dina = {96'd0, 16'd57081, 16'd46372, 16'd47067, 16'd65180, 16'd4126, 16'd17911, 16'd32010, 16'd2754, 16'd19472, 16'd54616}; // indx = 5101
    #10;
    addra = 32'd163264;
    dina = {96'd0, 16'd54749, 16'd40118, 16'd43139, 16'd13607, 16'd9063, 16'd22309, 16'd33829, 16'd25917, 16'd57444, 16'd62192}; // indx = 5102
    #10;
    addra = 32'd163296;
    dina = {96'd0, 16'd12789, 16'd48645, 16'd15572, 16'd62984, 16'd63225, 16'd63839, 16'd27433, 16'd52867, 16'd26228, 16'd21254}; // indx = 5103
    #10;
    addra = 32'd163328;
    dina = {96'd0, 16'd1374, 16'd20133, 16'd15935, 16'd27866, 16'd60993, 16'd45420, 16'd20767, 16'd57493, 16'd16276, 16'd42853}; // indx = 5104
    #10;
    addra = 32'd163360;
    dina = {96'd0, 16'd12565, 16'd3507, 16'd57996, 16'd59183, 16'd40092, 16'd31272, 16'd47790, 16'd27354, 16'd29974, 16'd32997}; // indx = 5105
    #10;
    addra = 32'd163392;
    dina = {96'd0, 16'd6576, 16'd49398, 16'd47216, 16'd62292, 16'd32591, 16'd52048, 16'd32263, 16'd62842, 16'd9759, 16'd47101}; // indx = 5106
    #10;
    addra = 32'd163424;
    dina = {96'd0, 16'd55681, 16'd27857, 16'd30867, 16'd3504, 16'd62414, 16'd7293, 16'd62670, 16'd43913, 16'd45418, 16'd4225}; // indx = 5107
    #10;
    addra = 32'd163456;
    dina = {96'd0, 16'd40533, 16'd30155, 16'd54820, 16'd58890, 16'd47818, 16'd34693, 16'd42329, 16'd5825, 16'd56970, 16'd4080}; // indx = 5108
    #10;
    addra = 32'd163488;
    dina = {96'd0, 16'd401, 16'd21849, 16'd3955, 16'd7214, 16'd6643, 16'd13217, 16'd3847, 16'd17356, 16'd9682, 16'd63441}; // indx = 5109
    #10;
    addra = 32'd163520;
    dina = {96'd0, 16'd17958, 16'd7091, 16'd19350, 16'd24295, 16'd39702, 16'd59264, 16'd10601, 16'd40776, 16'd29863, 16'd45586}; // indx = 5110
    #10;
    addra = 32'd163552;
    dina = {96'd0, 16'd44463, 16'd2226, 16'd59993, 16'd52812, 16'd17345, 16'd35821, 16'd465, 16'd39675, 16'd23300, 16'd17514}; // indx = 5111
    #10;
    addra = 32'd163584;
    dina = {96'd0, 16'd10544, 16'd55737, 16'd56824, 16'd9322, 16'd21999, 16'd52436, 16'd61651, 16'd36070, 16'd24064, 16'd54446}; // indx = 5112
    #10;
    addra = 32'd163616;
    dina = {96'd0, 16'd4658, 16'd18164, 16'd35611, 16'd45904, 16'd26062, 16'd25643, 16'd55976, 16'd14397, 16'd51191, 16'd2831}; // indx = 5113
    #10;
    addra = 32'd163648;
    dina = {96'd0, 16'd65311, 16'd4834, 16'd27465, 16'd55171, 16'd5423, 16'd10380, 16'd34792, 16'd63003, 16'd24191, 16'd62831}; // indx = 5114
    #10;
    addra = 32'd163680;
    dina = {96'd0, 16'd33236, 16'd3002, 16'd58922, 16'd33300, 16'd7968, 16'd45799, 16'd25951, 16'd29150, 16'd38760, 16'd5149}; // indx = 5115
    #10;
    addra = 32'd163712;
    dina = {96'd0, 16'd47634, 16'd26783, 16'd38517, 16'd15703, 16'd21694, 16'd37195, 16'd34991, 16'd65164, 16'd33428, 16'd12746}; // indx = 5116
    #10;
    addra = 32'd163744;
    dina = {96'd0, 16'd46171, 16'd44394, 16'd63722, 16'd22072, 16'd57849, 16'd21879, 16'd11744, 16'd61308, 16'd11146, 16'd34121}; // indx = 5117
    #10;
    addra = 32'd163776;
    dina = {96'd0, 16'd50938, 16'd35977, 16'd35043, 16'd26658, 16'd44129, 16'd44920, 16'd53235, 16'd38980, 16'd50175, 16'd24115}; // indx = 5118
    #10;
    addra = 32'd163808;
    dina = {96'd0, 16'd58834, 16'd58834, 16'd13271, 16'd3328, 16'd43408, 16'd11781, 16'd54877, 16'd45802, 16'd31296, 16'd12654}; // indx = 5119
    #10;

    ena = 0;
    wea = 0;

    #50;
    start = 1;
    #10;
    start = 0;

    #500000 $finish;
  end

  always #5 clk = ~clk;

endmodule
