`timescale 1ns / 1ps

module margin_sampling10(
  input  wire clk,
  input  wire rst_n,
  // *** CONTROL AND STATUS PORT ***
  output wire ready,
  input  wire start,
  // *** DATA INPUT PORT ***
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA CLK" *)  output wire clka,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA RST" *)  output wire rsta,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA EN" *)   output wire ena,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA ADDR" *) output wire [31:0] addra,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA DIN" *)  output wire [255:0] dina,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA WE" *)   output wire [31:0] wea,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA DOUT" *) input  wire [255:0] douta,
  // *** DATA OUTPUT PORT ***
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB CLK" *)  output wire clkb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB RST" *)  output wire rstb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB EN" *)   output wire enb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB ADDR" *) output wire [31:0] addrb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB DIN" *)  output wire [31:0] dinb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB WE" *)   output wire [3:0] web,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB DOUT" *) input  wire [31:0] doutb
);
  
  //local parameters
  localparam DATA_WIDTH = 16;
  localparam BATCH_SIZE = 1024;
  localparam MAX_DATA_LENGTH = 10*BATCH_SIZE;
  localparam DATA_LENGTH = 10240;
  localparam ADDR_WIDTH_PORTA = 32;
  localparam ADDR_INCR_PORTA = 32;
  localparam ADDR_WIDTH_PORTB = 32;
  localparam ADDR_INCR_PORTB = 4;
  localparam N_REGISTERS = 128;
  localparam N_REGISTERSBANKS = 8;
  localparam INDX_WIDTH = $clog2(MAX_DATA_LENGTH);
  localparam ADDR_WIDTH = $clog2(N_REGISTERS);
  localparam MARGIN_PIPELINE_DEPTH = 7;
  
  //wires
  wire startrising;
  
  wire [DATA_WIDTH-1:0] din0, din1, din2, din3, din4, din5, din6, din7, din8, din9;
  wire [DATA_WIDTH-1:0] rdin0, rdin1, rdin2, rdin3, rdin4, rdin5, rdin6, rdin7, rdin8, rdin9;
  wire [DATA_WIDTH-1:0] mrgn;
  
  wire trigmax;
  wire enaw;
  wire [31:0] weaw;
  wire enbw;
  wire [3:0] webw;
  wire cntaddraen;
  wire mrgnpipelineen;
  wire cntindxen;  
  wire cntren;
  wire cntrben;
  wire rsrc;  
  wire rbsrc;
  wire decrsrc;
  wire mrgnsrc; 
  wire trigmtree;
  wire cntouten;
  wire cntaddrben;
  
  wire [ADDR_WIDTH_PORTA-1:0] addraw;
  wire [ADDR_WIDTH_PORTB-1:0] addrbw;
  wire [INDX_WIDTH-1:0] mrgnindx;
  wire [INDX_WIDTH-1:0] indx;
  wire [$clog2(N_REGISTERS)-1:0] cntr;
  wire [$clog2(N_REGISTERSBANKS)-1:0] cntrb;
  wire [$clog2(N_REGISTERS)-1:0] decrsrcmuxout;
  wire [N_REGISTERS-1:0] decr;
  wire [N_REGISTERSBANKS-1:0] decrb;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] mrgnsrcmuxout;
  wire [N_REGISTERS-1:0] rsrcmuxout;
  wire [N_REGISTERSBANKS-1:0] rbsrcmuxout;
  
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] r0tomtree0, r1tomtree0, r2tomtree0, r3tomtree0, r4tomtree0, r5tomtree0,
  r6tomtree0, r7tomtree0, r8tomtree0, r9tomtree0, r10tomtree0, r11tomtree0, r12tomtree0, r13tomtree0, r14tomtree0, r15tomtree0,
  r16tomtree0, r17tomtree0, r18tomtree0, r19tomtree0, r20tomtree0, r21tomtree0, r22tomtree0, r23tomtree0, r24tomtree0, r25tomtree0,
  r26tomtree0, r27tomtree0, r28tomtree0, r29tomtree0, r30tomtree0, r31tomtree0, r32tomtree0, r33tomtree0, r34tomtree0, r35tomtree0,
  r36tomtree0, r37tomtree0, r38tomtree0, r39tomtree0, r40tomtree0, r41tomtree0, r42tomtree0, r43tomtree0, r44tomtree0, r45tomtree0,
  r46tomtree0, r47tomtree0, r48tomtree0, r49tomtree0, r50tomtree0, r51tomtree0, r52tomtree0, r53tomtree0, r54tomtree0, r55tomtree0,
  r56tomtree0, r57tomtree0, r58tomtree0, r59tomtree0, r60tomtree0, r61tomtree0, r62tomtree0, r63tomtree0, r64tomtree0, r65tomtree0,
  r66tomtree0, r67tomtree0, r68tomtree0, r69tomtree0, r70tomtree0, r71tomtree0, r72tomtree0, r73tomtree0, r74tomtree0, r75tomtree0,
  r76tomtree0, r77tomtree0, r78tomtree0, r79tomtree0, r80tomtree0, r81tomtree0, r82tomtree0, r83tomtree0, r84tomtree0, r85tomtree0,
  r86tomtree0, r87tomtree0, r88tomtree0, r89tomtree0, r90tomtree0, r91tomtree0, r92tomtree0, r93tomtree0, r94tomtree0, r95tomtree0,
  r96tomtree0, r97tomtree0, r98tomtree0, r99tomtree0, r100tomtree0, r101tomtree0, r102tomtree0, r103tomtree0, r104tomtree0, r105tomtree0,
  r106tomtree0, r107tomtree0, r108tomtree0, r109tomtree0, r110tomtree0, r111tomtree0, r112tomtree0, r113tomtree0, r114tomtree0, r115tomtree0,
  r116tomtree0, r117tomtree0, r118tomtree0, r119tomtree0, r120tomtree0, r121tomtree0, r122tomtree0, r123tomtree0, r124tomtree0, r125tomtree0,
  r126tomtree0, r127tomtree0, r128tomtree1, r129tomtree1, r130tomtree1, r131tomtree1, r132tomtree1, r133tomtree1, r134tomtree1, r135tomtree1,
  r136tomtree1, r137tomtree1, r138tomtree1, r139tomtree1, r140tomtree1, r141tomtree1, r142tomtree1, r143tomtree1, r144tomtree1, r145tomtree1,
  r146tomtree1, r147tomtree1, r148tomtree1, r149tomtree1, r150tomtree1, r151tomtree1, r152tomtree1, r153tomtree1, r154tomtree1, r155tomtree1,
  r156tomtree1, r157tomtree1, r158tomtree1, r159tomtree1, r160tomtree1, r161tomtree1, r162tomtree1, r163tomtree1, r164tomtree1, r165tomtree1,
  r166tomtree1, r167tomtree1, r168tomtree1, r169tomtree1, r170tomtree1, r171tomtree1, r172tomtree1, r173tomtree1, r174tomtree1, r175tomtree1,
  r176tomtree1, r177tomtree1, r178tomtree1, r179tomtree1, r180tomtree1, r181tomtree1, r182tomtree1, r183tomtree1, r184tomtree1, r185tomtree1,
  r186tomtree1, r187tomtree1, r188tomtree1, r189tomtree1, r190tomtree1, r191tomtree1, r192tomtree1, r193tomtree1, r194tomtree1, r195tomtree1,
  r196tomtree1, r197tomtree1, r198tomtree1, r199tomtree1, r200tomtree1, r201tomtree1, r202tomtree1, r203tomtree1, r204tomtree1, r205tomtree1,
  r206tomtree1, r207tomtree1, r208tomtree1, r209tomtree1, r210tomtree1, r211tomtree1, r212tomtree1, r213tomtree1, r214tomtree1, r215tomtree1,
  r216tomtree1, r217tomtree1, r218tomtree1, r219tomtree1, r220tomtree1, r221tomtree1, r222tomtree1, r223tomtree1, r224tomtree1, r225tomtree1,
  r226tomtree1, r227tomtree1, r228tomtree1, r229tomtree1, r230tomtree1, r231tomtree1, r232tomtree1, r233tomtree1, r234tomtree1, r235tomtree1,
  r236tomtree1, r237tomtree1, r238tomtree1, r239tomtree1, r240tomtree1, r241tomtree1, r242tomtree1, r243tomtree1, r244tomtree1, r245tomtree1,
  r246tomtree1, r247tomtree1, r248tomtree1, r249tomtree1, r250tomtree1, r251tomtree1, r252tomtree1, r253tomtree1, r254tomtree1, r255tomtree1,
  r256tomtree2, r257tomtree2, r258tomtree2, r259tomtree2, r260tomtree2, r261tomtree2, r262tomtree2, r263tomtree2, r264tomtree2, r265tomtree2,
  r266tomtree2, r267tomtree2, r268tomtree2, r269tomtree2, r270tomtree2, r271tomtree2, r272tomtree2, r273tomtree2, r274tomtree2, r275tomtree2,
  r276tomtree2, r277tomtree2, r278tomtree2, r279tomtree2, r280tomtree2, r281tomtree2, r282tomtree2, r283tomtree2, r284tomtree2, r285tomtree2,
  r286tomtree2, r287tomtree2, r288tomtree2, r289tomtree2, r290tomtree2, r291tomtree2, r292tomtree2, r293tomtree2, r294tomtree2, r295tomtree2,
  r296tomtree2, r297tomtree2, r298tomtree2, r299tomtree2, r300tomtree2, r301tomtree2, r302tomtree2, r303tomtree2, r304tomtree2, r305tomtree2,
  r306tomtree2, r307tomtree2, r308tomtree2, r309tomtree2, r310tomtree2, r311tomtree2, r312tomtree2, r313tomtree2, r314tomtree2, r315tomtree2,
  r316tomtree2, r317tomtree2, r318tomtree2, r319tomtree2, r320tomtree2, r321tomtree2, r322tomtree2, r323tomtree2, r324tomtree2, r325tomtree2,
  r326tomtree2, r327tomtree2, r328tomtree2, r329tomtree2, r330tomtree2, r331tomtree2, r332tomtree2, r333tomtree2, r334tomtree2, r335tomtree2,
  r336tomtree2, r337tomtree2, r338tomtree2, r339tomtree2, r340tomtree2, r341tomtree2, r342tomtree2, r343tomtree2, r344tomtree2, r345tomtree2,
  r346tomtree2, r347tomtree2, r348tomtree2, r349tomtree2, r350tomtree2, r351tomtree2, r352tomtree2, r353tomtree2, r354tomtree2, r355tomtree2,
  r356tomtree2, r357tomtree2, r358tomtree2, r359tomtree2, r360tomtree2, r361tomtree2, r362tomtree2, r363tomtree2, r364tomtree2, r365tomtree2,
  r366tomtree2, r367tomtree2, r368tomtree2, r369tomtree2, r370tomtree2, r371tomtree2, r372tomtree2, r373tomtree2, r374tomtree2, r375tomtree2,
  r376tomtree2, r377tomtree2, r378tomtree2, r379tomtree2, r380tomtree2, r381tomtree2, r382tomtree2, r383tomtree2, r384tomtree3, r385tomtree3,
  r386tomtree3, r387tomtree3, r388tomtree3, r389tomtree3, r390tomtree3, r391tomtree3, r392tomtree3, r393tomtree3, r394tomtree3, r395tomtree3,
  r396tomtree3, r397tomtree3, r398tomtree3, r399tomtree3, r400tomtree3, r401tomtree3, r402tomtree3, r403tomtree3, r404tomtree3, r405tomtree3,
  r406tomtree3, r407tomtree3, r408tomtree3, r409tomtree3, r410tomtree3, r411tomtree3, r412tomtree3, r413tomtree3, r414tomtree3, r415tomtree3,
  r416tomtree3, r417tomtree3, r418tomtree3, r419tomtree3, r420tomtree3, r421tomtree3, r422tomtree3, r423tomtree3, r424tomtree3, r425tomtree3,
  r426tomtree3, r427tomtree3, r428tomtree3, r429tomtree3, r430tomtree3, r431tomtree3, r432tomtree3, r433tomtree3, r434tomtree3, r435tomtree3,
  r436tomtree3, r437tomtree3, r438tomtree3, r439tomtree3, r440tomtree3, r441tomtree3, r442tomtree3, r443tomtree3, r444tomtree3, r445tomtree3,
  r446tomtree3, r447tomtree3, r448tomtree3, r449tomtree3, r450tomtree3, r451tomtree3, r452tomtree3, r453tomtree3, r454tomtree3, r455tomtree3,
  r456tomtree3, r457tomtree3, r458tomtree3, r459tomtree3, r460tomtree3, r461tomtree3, r462tomtree3, r463tomtree3, r464tomtree3, r465tomtree3,
  r466tomtree3, r467tomtree3, r468tomtree3, r469tomtree3, r470tomtree3, r471tomtree3, r472tomtree3, r473tomtree3, r474tomtree3, r475tomtree3,
  r476tomtree3, r477tomtree3, r478tomtree3, r479tomtree3, r480tomtree3, r481tomtree3, r482tomtree3, r483tomtree3, r484tomtree3, r485tomtree3,
  r486tomtree3, r487tomtree3, r488tomtree3, r489tomtree3, r490tomtree3, r491tomtree3, r492tomtree3, r493tomtree3, r494tomtree3, r495tomtree3,
  r496tomtree3, r497tomtree3, r498tomtree3, r499tomtree3, r500tomtree3, r501tomtree3, r502tomtree3, r503tomtree3, r504tomtree3, r505tomtree3,
  r506tomtree3, r507tomtree3, r508tomtree3, r509tomtree3, r510tomtree3, r511tomtree3, r512tomtree4, r513tomtree4, r514tomtree4, r515tomtree4,
  r516tomtree4, r517tomtree4, r518tomtree4, r519tomtree4, r520tomtree4, r521tomtree4, r522tomtree4, r523tomtree4, r524tomtree4, r525tomtree4,
  r526tomtree4, r527tomtree4, r528tomtree4, r529tomtree4, r530tomtree4, r531tomtree4, r532tomtree4, r533tomtree4, r534tomtree4, r535tomtree4,
  r536tomtree4, r537tomtree4, r538tomtree4, r539tomtree4, r540tomtree4, r541tomtree4, r542tomtree4, r543tomtree4, r544tomtree4, r545tomtree4,
  r546tomtree4, r547tomtree4, r548tomtree4, r549tomtree4, r550tomtree4, r551tomtree4, r552tomtree4, r553tomtree4, r554tomtree4, r555tomtree4,
  r556tomtree4, r557tomtree4, r558tomtree4, r559tomtree4, r560tomtree4, r561tomtree4, r562tomtree4, r563tomtree4, r564tomtree4, r565tomtree4,
  r566tomtree4, r567tomtree4, r568tomtree4, r569tomtree4, r570tomtree4, r571tomtree4, r572tomtree4, r573tomtree4, r574tomtree4, r575tomtree4,
  r576tomtree4, r577tomtree4, r578tomtree4, r579tomtree4, r580tomtree4, r581tomtree4, r582tomtree4, r583tomtree4, r584tomtree4, r585tomtree4,
  r586tomtree4, r587tomtree4, r588tomtree4, r589tomtree4, r590tomtree4, r591tomtree4, r592tomtree4, r593tomtree4, r594tomtree4, r595tomtree4,
  r596tomtree4, r597tomtree4, r598tomtree4, r599tomtree4, r600tomtree4, r601tomtree4, r602tomtree4, r603tomtree4, r604tomtree4, r605tomtree4,
  r606tomtree4, r607tomtree4, r608tomtree4, r609tomtree4, r610tomtree4, r611tomtree4, r612tomtree4, r613tomtree4, r614tomtree4, r615tomtree4,
  r616tomtree4, r617tomtree4, r618tomtree4, r619tomtree4, r620tomtree4, r621tomtree4, r622tomtree4, r623tomtree4, r624tomtree4, r625tomtree4,
  r626tomtree4, r627tomtree4, r628tomtree4, r629tomtree4, r630tomtree4, r631tomtree4, r632tomtree4, r633tomtree4, r634tomtree4, r635tomtree4,
  r636tomtree4, r637tomtree4, r638tomtree4, r639tomtree4, r640tomtree5, r641tomtree5, r642tomtree5, r643tomtree5, r644tomtree5, r645tomtree5,
  r646tomtree5, r647tomtree5, r648tomtree5, r649tomtree5, r650tomtree5, r651tomtree5, r652tomtree5, r653tomtree5, r654tomtree5, r655tomtree5,
  r656tomtree5, r657tomtree5, r658tomtree5, r659tomtree5, r660tomtree5, r661tomtree5, r662tomtree5, r663tomtree5, r664tomtree5, r665tomtree5,
  r666tomtree5, r667tomtree5, r668tomtree5, r669tomtree5, r670tomtree5, r671tomtree5, r672tomtree5, r673tomtree5, r674tomtree5, r675tomtree5,
  r676tomtree5, r677tomtree5, r678tomtree5, r679tomtree5, r680tomtree5, r681tomtree5, r682tomtree5, r683tomtree5, r684tomtree5, r685tomtree5,
  r686tomtree5, r687tomtree5, r688tomtree5, r689tomtree5, r690tomtree5, r691tomtree5, r692tomtree5, r693tomtree5, r694tomtree5, r695tomtree5,
  r696tomtree5, r697tomtree5, r698tomtree5, r699tomtree5, r700tomtree5, r701tomtree5, r702tomtree5, r703tomtree5, r704tomtree5, r705tomtree5,
  r706tomtree5, r707tomtree5, r708tomtree5, r709tomtree5, r710tomtree5, r711tomtree5, r712tomtree5, r713tomtree5, r714tomtree5, r715tomtree5,
  r716tomtree5, r717tomtree5, r718tomtree5, r719tomtree5, r720tomtree5, r721tomtree5, r722tomtree5, r723tomtree5, r724tomtree5, r725tomtree5,
  r726tomtree5, r727tomtree5, r728tomtree5, r729tomtree5, r730tomtree5, r731tomtree5, r732tomtree5, r733tomtree5, r734tomtree5, r735tomtree5,
  r736tomtree5, r737tomtree5, r738tomtree5, r739tomtree5, r740tomtree5, r741tomtree5, r742tomtree5, r743tomtree5, r744tomtree5, r745tomtree5,
  r746tomtree5, r747tomtree5, r748tomtree5, r749tomtree5, r750tomtree5, r751tomtree5, r752tomtree5, r753tomtree5, r754tomtree5, r755tomtree5,
  r756tomtree5, r757tomtree5, r758tomtree5, r759tomtree5, r760tomtree5, r761tomtree5, r762tomtree5, r763tomtree5, r764tomtree5, r765tomtree5,
  r766tomtree5, r767tomtree5, r768tomtree6, r769tomtree6, r770tomtree6, r771tomtree6, r772tomtree6, r773tomtree6, r774tomtree6, r775tomtree6,
  r776tomtree6, r777tomtree6, r778tomtree6, r779tomtree6, r780tomtree6, r781tomtree6, r782tomtree6, r783tomtree6, r784tomtree6, r785tomtree6,
  r786tomtree6, r787tomtree6, r788tomtree6, r789tomtree6, r790tomtree6, r791tomtree6, r792tomtree6, r793tomtree6, r794tomtree6, r795tomtree6,
  r796tomtree6, r797tomtree6, r798tomtree6, r799tomtree6, r800tomtree6, r801tomtree6, r802tomtree6, r803tomtree6, r804tomtree6, r805tomtree6,
  r806tomtree6, r807tomtree6, r808tomtree6, r809tomtree6, r810tomtree6, r811tomtree6, r812tomtree6, r813tomtree6, r814tomtree6, r815tomtree6,
  r816tomtree6, r817tomtree6, r818tomtree6, r819tomtree6, r820tomtree6, r821tomtree6, r822tomtree6, r823tomtree6, r824tomtree6, r825tomtree6,
  r826tomtree6, r827tomtree6, r828tomtree6, r829tomtree6, r830tomtree6, r831tomtree6, r832tomtree6, r833tomtree6, r834tomtree6, r835tomtree6,
  r836tomtree6, r837tomtree6, r838tomtree6, r839tomtree6, r840tomtree6, r841tomtree6, r842tomtree6, r843tomtree6, r844tomtree6, r845tomtree6,
  r846tomtree6, r847tomtree6, r848tomtree6, r849tomtree6, r850tomtree6, r851tomtree6, r852tomtree6, r853tomtree6, r854tomtree6, r855tomtree6,
  r856tomtree6, r857tomtree6, r858tomtree6, r859tomtree6, r860tomtree6, r861tomtree6, r862tomtree6, r863tomtree6, r864tomtree6, r865tomtree6,
  r866tomtree6, r867tomtree6, r868tomtree6, r869tomtree6, r870tomtree6, r871tomtree6, r872tomtree6, r873tomtree6, r874tomtree6, r875tomtree6,
  r876tomtree6, r877tomtree6, r878tomtree6, r879tomtree6, r880tomtree6, r881tomtree6, r882tomtree6, r883tomtree6, r884tomtree6, r885tomtree6,
  r886tomtree6, r887tomtree6, r888tomtree6, r889tomtree6, r890tomtree6, r891tomtree6, r892tomtree6, r893tomtree6, r894tomtree6, r895tomtree6,
  r896tomtree7, r897tomtree7, r898tomtree7, r899tomtree7, r900tomtree7, r901tomtree7, r902tomtree7, r903tomtree7, r904tomtree7, r905tomtree7,
  r906tomtree7, r907tomtree7, r908tomtree7, r909tomtree7, r910tomtree7, r911tomtree7, r912tomtree7, r913tomtree7, r914tomtree7, r915tomtree7,
  r916tomtree7, r917tomtree7, r918tomtree7, r919tomtree7, r920tomtree7, r921tomtree7, r922tomtree7, r923tomtree7, r924tomtree7, r925tomtree7,
  r926tomtree7, r927tomtree7, r928tomtree7, r929tomtree7, r930tomtree7, r931tomtree7, r932tomtree7, r933tomtree7, r934tomtree7, r935tomtree7,
  r936tomtree7, r937tomtree7, r938tomtree7, r939tomtree7, r940tomtree7, r941tomtree7, r942tomtree7, r943tomtree7, r944tomtree7, r945tomtree7,
  r946tomtree7, r947tomtree7, r948tomtree7, r949tomtree7, r950tomtree7, r951tomtree7, r952tomtree7, r953tomtree7, r954tomtree7, r955tomtree7,
  r956tomtree7, r957tomtree7, r958tomtree7, r959tomtree7, r960tomtree7, r961tomtree7, r962tomtree7, r963tomtree7, r964tomtree7, r965tomtree7,
  r966tomtree7, r967tomtree7, r968tomtree7, r969tomtree7, r970tomtree7, r971tomtree7, r972tomtree7, r973tomtree7, r974tomtree7, r975tomtree7,
  r976tomtree7, r977tomtree7, r978tomtree7, r979tomtree7, r980tomtree7, r981tomtree7, r982tomtree7, r983tomtree7, r984tomtree7, r985tomtree7,
  r986tomtree7, r987tomtree7, r988tomtree7, r989tomtree7, r990tomtree7, r991tomtree7, r992tomtree7, r993tomtree7, r994tomtree7, r995tomtree7,
  r996tomtree7, r997tomtree7, r998tomtree7, r999tomtree7, r1000tomtree7, r1001tomtree7, r1002tomtree7, r1003tomtree7, r1004tomtree7, r1005tomtree7,
  r1006tomtree7, r1007tomtree7, r1008tomtree7, r1009tomtree7, r1010tomtree7, r1011tomtree7, r1012tomtree7, r1013tomtree7, r1014tomtree7, r1015tomtree7,
  r1016tomtree7, r1017tomtree7, r1018tomtree7, r1019tomtree7, r1020tomtree7, r1021tomtree7, r1022tomtree7, r1023tomtree7;
  
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] mtree0tomaxsrcmux, mtree1tomaxsrcmux, mtree2tomaxsrcmux, 
  mtree3tomaxsrcmux, mtree4tomaxsrcmux, mtree5tomaxsrcmux, mtree6tomaxsrcmux, mtree7tomaxsrcmux;
  
  wire [N_REGISTERSBANKS-1:0] trigmtreesrcmuxout;
  wire [N_REGISTERSBANKS-1:0] trigmtreeold;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] maxsrcmuxtocmp;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] mrgncmp;
  wire [$clog2(N_REGISTERS)-1:0] rcmp; 
  wire [$clog2(BATCH_SIZE)-1:0] cntout;
  
  //start rising
  reg startold;
  always @(posedge clk) begin
    startold <= start;
  end
  assign startrising = !startold && start;
  
  controller #(.DATA_LENGTH(DATA_LENGTH), .MARGIN_PIPELINE_DEPTH(MARGIN_PIPELINE_DEPTH), .N_REGISTERS(N_REGISTERS), .BATCH_SIZE(BATCH_SIZE), .N_REGISTERSBANKS(N_REGISTERSBANKS)) Cntr(
    .clk(clk),
    .rst_n(rst_n),
    .Start(startrising),
    .MTreeSrc(trigmax),
    .Ready(ready),
    .EnA(enaw),
    .WeA(weaw),
    .EnB(enbw),
    .WeB(webw),
    .CntAddrAEn(cntaddraen),
    .MrgnPipelineEn(mrgnpipelineen),
    .CntIndxEn(cntindxen),
    .CntREn(cntren),
    .CntRBEn(cntrben),
    .RSrc(rsrc),
    .RBSrc(rbsrc),
    .DecRSrc(decrsrc),
    .MrgnSrc(mrgnsrc),
    .TrigMTree(trigmtree),
    .CntOutEn(cntouten),
    .CntAddrBEn(cntaddrben)
  );

  //bram input port
  assign clka = clk;
  assign rsta = ~rst_n;
  assign ena = enaw;
  assign addra = addraw;
  assign dina = 0;
  assign wea = weaw;
  
  counter_addr #(.INCR(ADDR_INCR_PORTA), .ADDR_WIDTH(ADDR_WIDTH_PORTA)) CntAddrA(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntaddraen),
    .cnt(addraw)
  );
  
  assign din0 = douta[15:0];
  assign din1 = douta[31:16];
  assign din2 = douta[47:32];
  assign din3 = douta[63:48];
  assign din4 = douta[79:64];
  assign din5 = douta[95:80];
  assign din6 = douta[111:96];
  assign din7 = douta[127:112];
  assign din8 = douta[143:128];
  assign din9 = douta[159:144];
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn0(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din0),
    .dout(rdin0)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn1(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din1),
    .dout(rdin1)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn2(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din2),
    .dout(rdin2)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn3(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din3),
    .dout(rdin3)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn4(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din4),
    .dout(rdin4)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn5(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din5),
    .dout(rdin5)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn6(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din6),
    .dout(rdin6)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn7(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din7),
    .dout(rdin7)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn8(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din8),
    .dout(rdin8)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn9(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din9),
    .dout(rdin9)
  );
  
  margin_pipeline10 #(.DATA_WIDTH(DATA_WIDTH)) MrgnPipeline(
    .clk(clk),
    .rst_n(rst_n),
    .en(mrgnpipelineen),
    .din0(rdin0),
    .din1(rdin1),
    .din2(rdin2),
    .din3(rdin3),
    .din4(rdin4),
    .din5(rdin5),
    .din6(rdin6),
    .din7(rdin7),
    .din8(rdin8),
    .din9(rdin9),
    .margin(mrgn)
  );
  
  counter_indx #(.INCR(1), .CNT_WIDTH(INDX_WIDTH)) CntIndx(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntindxen),
    .cnt(mrgnindx)
  );
  
  counter_r #(.MAX_CNT(N_REGISTERS), .INCR(1), .N_REGISTERSBANKS(N_REGISTERSBANKS)) CntR(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntren),
    .cnt(cntr)
  );

  mux2 #(.DATA_WIDTH($clog2(N_REGISTERS))) DecRSrcMux(
    .din0(cntr), 
    .din1(rcmp), 
    .sel(decrsrc), 
    .dout(decrsrcmuxout)
  );

  decoder #(.IN_WIDTH($clog2(N_REGISTERS))) DecR(
    .din(decrsrcmuxout), 
    .dout(decr)
  );

  counter_rb #(.MAX_CNT(N_REGISTERSBANKS), .INCR(1)) CntRB(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntrben),
    .cnt(cntrb)
  );

  decoder #(.IN_WIDTH($clog2(N_REGISTERSBANKS))) DecRB(
    .din(cntrb), 
    .dout(decrb)
  );

  mux2 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) MrgnSrcMux(
    .din0(mrgncmp), 
    .din1({cntr,mrgnindx,mrgn}), 
    .sel(!mrgnsrc), 
    .dout(mrgnsrcmuxout)
  );

  mux2 #(.DATA_WIDTH(N_REGISTERS)) RSrcMux(
    .din0('b0), 
    .din1(decr), 
    .sel(rsrc), 
    .dout(rsrcmuxout)
  );

  mux2 #(.DATA_WIDTH(N_REGISTERSBANKS)) RBSrcMux(
    .din0('b0), 
    .din1(decrb), 
    .sel(rsrc), 
    .dout(rbsrcmuxout)
  );
  
  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_0(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[0]),
    .din(mrgnsrcmuxout),
    .dout0(r0tomtree0),
    .dout1(r1tomtree0),
    .dout2(r2tomtree0),
    .dout3(r3tomtree0),
    .dout4(r4tomtree0),
    .dout5(r5tomtree0),
    .dout6(r6tomtree0),
    .dout7(r7tomtree0),
    .dout8(r8tomtree0),
    .dout9(r9tomtree0),
    .dout10(r10tomtree0),
    .dout11(r11tomtree0),
    .dout12(r12tomtree0),
    .dout13(r13tomtree0),
    .dout14(r14tomtree0),
    .dout15(r15tomtree0),
    .dout16(r16tomtree0),
    .dout17(r17tomtree0),
    .dout18(r18tomtree0),
    .dout19(r19tomtree0),
    .dout20(r20tomtree0),
    .dout21(r21tomtree0),
    .dout22(r22tomtree0),
    .dout23(r23tomtree0),
    .dout24(r24tomtree0),
    .dout25(r25tomtree0),
    .dout26(r26tomtree0),
    .dout27(r27tomtree0),
    .dout28(r28tomtree0),
    .dout29(r29tomtree0),
    .dout30(r30tomtree0),
    .dout31(r31tomtree0),
    .dout32(r32tomtree0),
    .dout33(r33tomtree0),
    .dout34(r34tomtree0),
    .dout35(r35tomtree0),
    .dout36(r36tomtree0),
    .dout37(r37tomtree0),
    .dout38(r38tomtree0),
    .dout39(r39tomtree0),
    .dout40(r40tomtree0),
    .dout41(r41tomtree0),
    .dout42(r42tomtree0),
    .dout43(r43tomtree0),
    .dout44(r44tomtree0),
    .dout45(r45tomtree0),
    .dout46(r46tomtree0),
    .dout47(r47tomtree0),
    .dout48(r48tomtree0),
    .dout49(r49tomtree0),
    .dout50(r50tomtree0),
    .dout51(r51tomtree0),
    .dout52(r52tomtree0),
    .dout53(r53tomtree0),
    .dout54(r54tomtree0),
    .dout55(r55tomtree0),
    .dout56(r56tomtree0),
    .dout57(r57tomtree0),
    .dout58(r58tomtree0),
    .dout59(r59tomtree0),
    .dout60(r60tomtree0),
    .dout61(r61tomtree0),
    .dout62(r62tomtree0),
    .dout63(r63tomtree0),
    .dout64(r64tomtree0),
    .dout65(r65tomtree0),
    .dout66(r66tomtree0),
    .dout67(r67tomtree0),
    .dout68(r68tomtree0),
    .dout69(r69tomtree0),
    .dout70(r70tomtree0),
    .dout71(r71tomtree0),
    .dout72(r72tomtree0),
    .dout73(r73tomtree0),
    .dout74(r74tomtree0),
    .dout75(r75tomtree0),
    .dout76(r76tomtree0),
    .dout77(r77tomtree0),
    .dout78(r78tomtree0),
    .dout79(r79tomtree0),
    .dout80(r80tomtree0),
    .dout81(r81tomtree0),
    .dout82(r82tomtree0),
    .dout83(r83tomtree0),
    .dout84(r84tomtree0),
    .dout85(r85tomtree0),
    .dout86(r86tomtree0),
    .dout87(r87tomtree0),
    .dout88(r88tomtree0),
    .dout89(r89tomtree0),
    .dout90(r90tomtree0),
    .dout91(r91tomtree0),
    .dout92(r92tomtree0),
    .dout93(r93tomtree0),
    .dout94(r94tomtree0),
    .dout95(r95tomtree0),
    .dout96(r96tomtree0),
    .dout97(r97tomtree0),
    .dout98(r98tomtree0),
    .dout99(r99tomtree0),
    .dout100(r100tomtree0),
    .dout101(r101tomtree0),
    .dout102(r102tomtree0),
    .dout103(r103tomtree0),
    .dout104(r104tomtree0),
    .dout105(r105tomtree0),
    .dout106(r106tomtree0),
    .dout107(r107tomtree0),
    .dout108(r108tomtree0),
    .dout109(r109tomtree0),
    .dout110(r110tomtree0),
    .dout111(r111tomtree0),
    .dout112(r112tomtree0),
    .dout113(r113tomtree0),
    .dout114(r114tomtree0),
    .dout115(r115tomtree0),
    .dout116(r116tomtree0),
    .dout117(r117tomtree0),
    .dout118(r118tomtree0),
    .dout119(r119tomtree0),
    .dout120(r120tomtree0),
    .dout121(r121tomtree0),
    .dout122(r122tomtree0),
    .dout123(r123tomtree0),
    .dout124(r124tomtree0),
    .dout125(r125tomtree0),
    .dout126(r126tomtree0),
    .dout127(r127tomtree0)
  );

  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_1(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[1]),
    .din(mrgnsrcmuxout),
    .dout0(r128tomtree1),
    .dout1(r129tomtree1),
    .dout2(r130tomtree1),
    .dout3(r131tomtree1),
    .dout4(r132tomtree1),
    .dout5(r133tomtree1),
    .dout6(r134tomtree1),
    .dout7(r135tomtree1),
    .dout8(r136tomtree1),
    .dout9(r137tomtree1),
    .dout10(r138tomtree1),
    .dout11(r139tomtree1),
    .dout12(r140tomtree1),
    .dout13(r141tomtree1),
    .dout14(r142tomtree1),
    .dout15(r143tomtree1),
    .dout16(r144tomtree1),
    .dout17(r145tomtree1),
    .dout18(r146tomtree1),
    .dout19(r147tomtree1),
    .dout20(r148tomtree1),
    .dout21(r149tomtree1),
    .dout22(r150tomtree1),
    .dout23(r151tomtree1),
    .dout24(r152tomtree1),
    .dout25(r153tomtree1),
    .dout26(r154tomtree1),
    .dout27(r155tomtree1),
    .dout28(r156tomtree1),
    .dout29(r157tomtree1),
    .dout30(r158tomtree1),
    .dout31(r159tomtree1),
    .dout32(r160tomtree1),
    .dout33(r161tomtree1),
    .dout34(r162tomtree1),
    .dout35(r163tomtree1),
    .dout36(r164tomtree1),
    .dout37(r165tomtree1),
    .dout38(r166tomtree1),
    .dout39(r167tomtree1),
    .dout40(r168tomtree1),
    .dout41(r169tomtree1),
    .dout42(r170tomtree1),
    .dout43(r171tomtree1),
    .dout44(r172tomtree1),
    .dout45(r173tomtree1),
    .dout46(r174tomtree1),
    .dout47(r175tomtree1),
    .dout48(r176tomtree1),
    .dout49(r177tomtree1),
    .dout50(r178tomtree1),
    .dout51(r179tomtree1),
    .dout52(r180tomtree1),
    .dout53(r181tomtree1),
    .dout54(r182tomtree1),
    .dout55(r183tomtree1),
    .dout56(r184tomtree1),
    .dout57(r185tomtree1),
    .dout58(r186tomtree1),
    .dout59(r187tomtree1),
    .dout60(r188tomtree1),
    .dout61(r189tomtree1),
    .dout62(r190tomtree1),
    .dout63(r191tomtree1),
    .dout64(r192tomtree1),
    .dout65(r193tomtree1),
    .dout66(r194tomtree1),
    .dout67(r195tomtree1),
    .dout68(r196tomtree1),
    .dout69(r197tomtree1),
    .dout70(r198tomtree1),
    .dout71(r199tomtree1),
    .dout72(r200tomtree1),
    .dout73(r201tomtree1),
    .dout74(r202tomtree1),
    .dout75(r203tomtree1),
    .dout76(r204tomtree1),
    .dout77(r205tomtree1),
    .dout78(r206tomtree1),
    .dout79(r207tomtree1),
    .dout80(r208tomtree1),
    .dout81(r209tomtree1),
    .dout82(r210tomtree1),
    .dout83(r211tomtree1),
    .dout84(r212tomtree1),
    .dout85(r213tomtree1),
    .dout86(r214tomtree1),
    .dout87(r215tomtree1),
    .dout88(r216tomtree1),
    .dout89(r217tomtree1),
    .dout90(r218tomtree1),
    .dout91(r219tomtree1),
    .dout92(r220tomtree1),
    .dout93(r221tomtree1),
    .dout94(r222tomtree1),
    .dout95(r223tomtree1),
    .dout96(r224tomtree1),
    .dout97(r225tomtree1),
    .dout98(r226tomtree1),
    .dout99(r227tomtree1),
    .dout100(r228tomtree1),
    .dout101(r229tomtree1),
    .dout102(r230tomtree1),
    .dout103(r231tomtree1),
    .dout104(r232tomtree1),
    .dout105(r233tomtree1),
    .dout106(r234tomtree1),
    .dout107(r235tomtree1),
    .dout108(r236tomtree1),
    .dout109(r237tomtree1),
    .dout110(r238tomtree1),
    .dout111(r239tomtree1),
    .dout112(r240tomtree1),
    .dout113(r241tomtree1),
    .dout114(r242tomtree1),
    .dout115(r243tomtree1),
    .dout116(r244tomtree1),
    .dout117(r245tomtree1),
    .dout118(r246tomtree1),
    .dout119(r247tomtree1),
    .dout120(r248tomtree1),
    .dout121(r249tomtree1),
    .dout122(r250tomtree1),
    .dout123(r251tomtree1),
    .dout124(r252tomtree1),
    .dout125(r253tomtree1),
    .dout126(r254tomtree1),
    .dout127(r255tomtree1)
  );

  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_2(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[2]),
    .din(mrgnsrcmuxout),
    .dout0(r256tomtree2),
    .dout1(r257tomtree2),
    .dout2(r258tomtree2),
    .dout3(r259tomtree2),
    .dout4(r260tomtree2),
    .dout5(r261tomtree2),
    .dout6(r262tomtree2),
    .dout7(r263tomtree2),
    .dout8(r264tomtree2),
    .dout9(r265tomtree2),
    .dout10(r266tomtree2),
    .dout11(r267tomtree2),
    .dout12(r268tomtree2),
    .dout13(r269tomtree2),
    .dout14(r270tomtree2),
    .dout15(r271tomtree2),
    .dout16(r272tomtree2),
    .dout17(r273tomtree2),
    .dout18(r274tomtree2),
    .dout19(r275tomtree2),
    .dout20(r276tomtree2),
    .dout21(r277tomtree2),
    .dout22(r278tomtree2),
    .dout23(r279tomtree2),
    .dout24(r280tomtree2),
    .dout25(r281tomtree2),
    .dout26(r282tomtree2),
    .dout27(r283tomtree2),
    .dout28(r284tomtree2),
    .dout29(r285tomtree2),
    .dout30(r286tomtree2),
    .dout31(r287tomtree2),
    .dout32(r288tomtree2),
    .dout33(r289tomtree2),
    .dout34(r290tomtree2),
    .dout35(r291tomtree2),
    .dout36(r292tomtree2),
    .dout37(r293tomtree2),
    .dout38(r294tomtree2),
    .dout39(r295tomtree2),
    .dout40(r296tomtree2),
    .dout41(r297tomtree2),
    .dout42(r298tomtree2),
    .dout43(r299tomtree2),
    .dout44(r300tomtree2),
    .dout45(r301tomtree2),
    .dout46(r302tomtree2),
    .dout47(r303tomtree2),
    .dout48(r304tomtree2),
    .dout49(r305tomtree2),
    .dout50(r306tomtree2),
    .dout51(r307tomtree2),
    .dout52(r308tomtree2),
    .dout53(r309tomtree2),
    .dout54(r310tomtree2),
    .dout55(r311tomtree2),
    .dout56(r312tomtree2),
    .dout57(r313tomtree2),
    .dout58(r314tomtree2),
    .dout59(r315tomtree2),
    .dout60(r316tomtree2),
    .dout61(r317tomtree2),
    .dout62(r318tomtree2),
    .dout63(r319tomtree2),
    .dout64(r320tomtree2),
    .dout65(r321tomtree2),
    .dout66(r322tomtree2),
    .dout67(r323tomtree2),
    .dout68(r324tomtree2),
    .dout69(r325tomtree2),
    .dout70(r326tomtree2),
    .dout71(r327tomtree2),
    .dout72(r328tomtree2),
    .dout73(r329tomtree2),
    .dout74(r330tomtree2),
    .dout75(r331tomtree2),
    .dout76(r332tomtree2),
    .dout77(r333tomtree2),
    .dout78(r334tomtree2),
    .dout79(r335tomtree2),
    .dout80(r336tomtree2),
    .dout81(r337tomtree2),
    .dout82(r338tomtree2),
    .dout83(r339tomtree2),
    .dout84(r340tomtree2),
    .dout85(r341tomtree2),
    .dout86(r342tomtree2),
    .dout87(r343tomtree2),
    .dout88(r344tomtree2),
    .dout89(r345tomtree2),
    .dout90(r346tomtree2),
    .dout91(r347tomtree2),
    .dout92(r348tomtree2),
    .dout93(r349tomtree2),
    .dout94(r350tomtree2),
    .dout95(r351tomtree2),
    .dout96(r352tomtree2),
    .dout97(r353tomtree2),
    .dout98(r354tomtree2),
    .dout99(r355tomtree2),
    .dout100(r356tomtree2),
    .dout101(r357tomtree2),
    .dout102(r358tomtree2),
    .dout103(r359tomtree2),
    .dout104(r360tomtree2),
    .dout105(r361tomtree2),
    .dout106(r362tomtree2),
    .dout107(r363tomtree2),
    .dout108(r364tomtree2),
    .dout109(r365tomtree2),
    .dout110(r366tomtree2),
    .dout111(r367tomtree2),
    .dout112(r368tomtree2),
    .dout113(r369tomtree2),
    .dout114(r370tomtree2),
    .dout115(r371tomtree2),
    .dout116(r372tomtree2),
    .dout117(r373tomtree2),
    .dout118(r374tomtree2),
    .dout119(r375tomtree2),
    .dout120(r376tomtree2),
    .dout121(r377tomtree2),
    .dout122(r378tomtree2),
    .dout123(r379tomtree2),
    .dout124(r380tomtree2),
    .dout125(r381tomtree2),
    .dout126(r382tomtree2),
    .dout127(r383tomtree2)
  );

  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_3(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[3]),
    .din(mrgnsrcmuxout),
    .dout0(r384tomtree3),
    .dout1(r385tomtree3),
    .dout2(r386tomtree3),
    .dout3(r387tomtree3),
    .dout4(r388tomtree3),
    .dout5(r389tomtree3),
    .dout6(r390tomtree3),
    .dout7(r391tomtree3),
    .dout8(r392tomtree3),
    .dout9(r393tomtree3),
    .dout10(r394tomtree3),
    .dout11(r395tomtree3),
    .dout12(r396tomtree3),
    .dout13(r397tomtree3),
    .dout14(r398tomtree3),
    .dout15(r399tomtree3),
    .dout16(r400tomtree3),
    .dout17(r401tomtree3),
    .dout18(r402tomtree3),
    .dout19(r403tomtree3),
    .dout20(r404tomtree3),
    .dout21(r405tomtree3),
    .dout22(r406tomtree3),
    .dout23(r407tomtree3),
    .dout24(r408tomtree3),
    .dout25(r409tomtree3),
    .dout26(r410tomtree3),
    .dout27(r411tomtree3),
    .dout28(r412tomtree3),
    .dout29(r413tomtree3),
    .dout30(r414tomtree3),
    .dout31(r415tomtree3),
    .dout32(r416tomtree3),
    .dout33(r417tomtree3),
    .dout34(r418tomtree3),
    .dout35(r419tomtree3),
    .dout36(r420tomtree3),
    .dout37(r421tomtree3),
    .dout38(r422tomtree3),
    .dout39(r423tomtree3),
    .dout40(r424tomtree3),
    .dout41(r425tomtree3),
    .dout42(r426tomtree3),
    .dout43(r427tomtree3),
    .dout44(r428tomtree3),
    .dout45(r429tomtree3),
    .dout46(r430tomtree3),
    .dout47(r431tomtree3),
    .dout48(r432tomtree3),
    .dout49(r433tomtree3),
    .dout50(r434tomtree3),
    .dout51(r435tomtree3),
    .dout52(r436tomtree3),
    .dout53(r437tomtree3),
    .dout54(r438tomtree3),
    .dout55(r439tomtree3),
    .dout56(r440tomtree3),
    .dout57(r441tomtree3),
    .dout58(r442tomtree3),
    .dout59(r443tomtree3),
    .dout60(r444tomtree3),
    .dout61(r445tomtree3),
    .dout62(r446tomtree3),
    .dout63(r447tomtree3),
    .dout64(r448tomtree3),
    .dout65(r449tomtree3),
    .dout66(r450tomtree3),
    .dout67(r451tomtree3),
    .dout68(r452tomtree3),
    .dout69(r453tomtree3),
    .dout70(r454tomtree3),
    .dout71(r455tomtree3),
    .dout72(r456tomtree3),
    .dout73(r457tomtree3),
    .dout74(r458tomtree3),
    .dout75(r459tomtree3),
    .dout76(r460tomtree3),
    .dout77(r461tomtree3),
    .dout78(r462tomtree3),
    .dout79(r463tomtree3),
    .dout80(r464tomtree3),
    .dout81(r465tomtree3),
    .dout82(r466tomtree3),
    .dout83(r467tomtree3),
    .dout84(r468tomtree3),
    .dout85(r469tomtree3),
    .dout86(r470tomtree3),
    .dout87(r471tomtree3),
    .dout88(r472tomtree3),
    .dout89(r473tomtree3),
    .dout90(r474tomtree3),
    .dout91(r475tomtree3),
    .dout92(r476tomtree3),
    .dout93(r477tomtree3),
    .dout94(r478tomtree3),
    .dout95(r479tomtree3),
    .dout96(r480tomtree3),
    .dout97(r481tomtree3),
    .dout98(r482tomtree3),
    .dout99(r483tomtree3),
    .dout100(r484tomtree3),
    .dout101(r485tomtree3),
    .dout102(r486tomtree3),
    .dout103(r487tomtree3),
    .dout104(r488tomtree3),
    .dout105(r489tomtree3),
    .dout106(r490tomtree3),
    .dout107(r491tomtree3),
    .dout108(r492tomtree3),
    .dout109(r493tomtree3),
    .dout110(r494tomtree3),
    .dout111(r495tomtree3),
    .dout112(r496tomtree3),
    .dout113(r497tomtree3),
    .dout114(r498tomtree3),
    .dout115(r499tomtree3),
    .dout116(r500tomtree3),
    .dout117(r501tomtree3),
    .dout118(r502tomtree3),
    .dout119(r503tomtree3),
    .dout120(r504tomtree3),
    .dout121(r505tomtree3),
    .dout122(r506tomtree3),
    .dout123(r507tomtree3),
    .dout124(r508tomtree3),
    .dout125(r509tomtree3),
    .dout126(r510tomtree3),
    .dout127(r511tomtree3)
  );
  
  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_4(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[4]),
    .din(mrgnsrcmuxout),
    .dout0(r512tomtree4),
    .dout1(r513tomtree4),
    .dout2(r514tomtree4),
    .dout3(r515tomtree4),
    .dout4(r516tomtree4),
    .dout5(r517tomtree4),
    .dout6(r518tomtree4),
    .dout7(r519tomtree4),
    .dout8(r520tomtree4),
    .dout9(r521tomtree4),
    .dout10(r522tomtree4),
    .dout11(r523tomtree4),
    .dout12(r524tomtree4),
    .dout13(r525tomtree4),
    .dout14(r526tomtree4),
    .dout15(r527tomtree4),
    .dout16(r528tomtree4),
    .dout17(r529tomtree4),
    .dout18(r530tomtree4),
    .dout19(r531tomtree4),
    .dout20(r532tomtree4),
    .dout21(r533tomtree4),
    .dout22(r534tomtree4),
    .dout23(r535tomtree4),
    .dout24(r536tomtree4),
    .dout25(r537tomtree4),
    .dout26(r538tomtree4),
    .dout27(r539tomtree4),
    .dout28(r540tomtree4),
    .dout29(r541tomtree4),
    .dout30(r542tomtree4),
    .dout31(r543tomtree4),
    .dout32(r544tomtree4),
    .dout33(r545tomtree4),
    .dout34(r546tomtree4),
    .dout35(r547tomtree4),
    .dout36(r548tomtree4),
    .dout37(r549tomtree4),
    .dout38(r550tomtree4),
    .dout39(r551tomtree4),
    .dout40(r552tomtree4),
    .dout41(r553tomtree4),
    .dout42(r554tomtree4),
    .dout43(r555tomtree4),
    .dout44(r556tomtree4),
    .dout45(r557tomtree4),
    .dout46(r558tomtree4),
    .dout47(r559tomtree4),
    .dout48(r560tomtree4),
    .dout49(r561tomtree4),
    .dout50(r562tomtree4),
    .dout51(r563tomtree4),
    .dout52(r564tomtree4),
    .dout53(r565tomtree4),
    .dout54(r566tomtree4),
    .dout55(r567tomtree4),
    .dout56(r568tomtree4),
    .dout57(r569tomtree4),
    .dout58(r570tomtree4),
    .dout59(r571tomtree4),
    .dout60(r572tomtree4),
    .dout61(r573tomtree4),
    .dout62(r574tomtree4),
    .dout63(r575tomtree4),
    .dout64(r576tomtree4),
    .dout65(r577tomtree4),
    .dout66(r578tomtree4),
    .dout67(r579tomtree4),
    .dout68(r580tomtree4),
    .dout69(r581tomtree4),
    .dout70(r582tomtree4),
    .dout71(r583tomtree4),
    .dout72(r584tomtree4),
    .dout73(r585tomtree4),
    .dout74(r586tomtree4),
    .dout75(r587tomtree4),
    .dout76(r588tomtree4),
    .dout77(r589tomtree4),
    .dout78(r590tomtree4),
    .dout79(r591tomtree4),
    .dout80(r592tomtree4),
    .dout81(r593tomtree4),
    .dout82(r594tomtree4),
    .dout83(r595tomtree4),
    .dout84(r596tomtree4),
    .dout85(r597tomtree4),
    .dout86(r598tomtree4),
    .dout87(r599tomtree4),
    .dout88(r600tomtree4),
    .dout89(r601tomtree4),
    .dout90(r602tomtree4),
    .dout91(r603tomtree4),
    .dout92(r604tomtree4),
    .dout93(r605tomtree4),
    .dout94(r606tomtree4),
    .dout95(r607tomtree4),
    .dout96(r608tomtree4),
    .dout97(r609tomtree4),
    .dout98(r610tomtree4),
    .dout99(r611tomtree4),
    .dout100(r612tomtree4),
    .dout101(r613tomtree4),
    .dout102(r614tomtree4),
    .dout103(r615tomtree4),
    .dout104(r616tomtree4),
    .dout105(r617tomtree4),
    .dout106(r618tomtree4),
    .dout107(r619tomtree4),
    .dout108(r620tomtree4),
    .dout109(r621tomtree4),
    .dout110(r622tomtree4),
    .dout111(r623tomtree4),
    .dout112(r624tomtree4),
    .dout113(r625tomtree4),
    .dout114(r626tomtree4),
    .dout115(r627tomtree4),
    .dout116(r628tomtree4),
    .dout117(r629tomtree4),
    .dout118(r630tomtree4),
    .dout119(r631tomtree4),
    .dout120(r632tomtree4),
    .dout121(r633tomtree4),
    .dout122(r634tomtree4),
    .dout123(r635tomtree4),
    .dout124(r636tomtree4),
    .dout125(r637tomtree4),
    .dout126(r638tomtree4),
    .dout127(r639tomtree4)
  );

  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_5(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[5]),
    .din(mrgnsrcmuxout),
    .dout0(r640tomtree5),
    .dout1(r641tomtree5),
    .dout2(r642tomtree5),
    .dout3(r643tomtree5),
    .dout4(r644tomtree5),
    .dout5(r645tomtree5),
    .dout6(r646tomtree5),
    .dout7(r647tomtree5),
    .dout8(r648tomtree5),
    .dout9(r649tomtree5),
    .dout10(r650tomtree5),
    .dout11(r651tomtree5),
    .dout12(r652tomtree5),
    .dout13(r653tomtree5),
    .dout14(r654tomtree5),
    .dout15(r655tomtree5),
    .dout16(r656tomtree5),
    .dout17(r657tomtree5),
    .dout18(r658tomtree5),
    .dout19(r659tomtree5),
    .dout20(r660tomtree5),
    .dout21(r661tomtree5),
    .dout22(r662tomtree5),
    .dout23(r663tomtree5),
    .dout24(r664tomtree5),
    .dout25(r665tomtree5),
    .dout26(r666tomtree5),
    .dout27(r667tomtree5),
    .dout28(r668tomtree5),
    .dout29(r669tomtree5),
    .dout30(r670tomtree5),
    .dout31(r671tomtree5),
    .dout32(r672tomtree5),
    .dout33(r673tomtree5),
    .dout34(r674tomtree5),
    .dout35(r675tomtree5),
    .dout36(r676tomtree5),
    .dout37(r677tomtree5),
    .dout38(r678tomtree5),
    .dout39(r679tomtree5),
    .dout40(r680tomtree5),
    .dout41(r681tomtree5),
    .dout42(r682tomtree5),
    .dout43(r683tomtree5),
    .dout44(r684tomtree5),
    .dout45(r685tomtree5),
    .dout46(r686tomtree5),
    .dout47(r687tomtree5),
    .dout48(r688tomtree5),
    .dout49(r689tomtree5),
    .dout50(r690tomtree5),
    .dout51(r691tomtree5),
    .dout52(r692tomtree5),
    .dout53(r693tomtree5),
    .dout54(r694tomtree5),
    .dout55(r695tomtree5),
    .dout56(r696tomtree5),
    .dout57(r697tomtree5),
    .dout58(r698tomtree5),
    .dout59(r699tomtree5),
    .dout60(r700tomtree5),
    .dout61(r701tomtree5),
    .dout62(r702tomtree5),
    .dout63(r703tomtree5),
    .dout64(r704tomtree5),
    .dout65(r705tomtree5),
    .dout66(r706tomtree5),
    .dout67(r707tomtree5),
    .dout68(r708tomtree5),
    .dout69(r709tomtree5),
    .dout70(r710tomtree5),
    .dout71(r711tomtree5),
    .dout72(r712tomtree5),
    .dout73(r713tomtree5),
    .dout74(r714tomtree5),
    .dout75(r715tomtree5),
    .dout76(r716tomtree5),
    .dout77(r717tomtree5),
    .dout78(r718tomtree5),
    .dout79(r719tomtree5),
    .dout80(r720tomtree5),
    .dout81(r721tomtree5),
    .dout82(r722tomtree5),
    .dout83(r723tomtree5),
    .dout84(r724tomtree5),
    .dout85(r725tomtree5),
    .dout86(r726tomtree5),
    .dout87(r727tomtree5),
    .dout88(r728tomtree5),
    .dout89(r729tomtree5),
    .dout90(r730tomtree5),
    .dout91(r731tomtree5),
    .dout92(r732tomtree5),
    .dout93(r733tomtree5),
    .dout94(r734tomtree5),
    .dout95(r735tomtree5),
    .dout96(r736tomtree5),
    .dout97(r737tomtree5),
    .dout98(r738tomtree5),
    .dout99(r739tomtree5),
    .dout100(r740tomtree5),
    .dout101(r741tomtree5),
    .dout102(r742tomtree5),
    .dout103(r743tomtree5),
    .dout104(r744tomtree5),
    .dout105(r745tomtree5),
    .dout106(r746tomtree5),
    .dout107(r747tomtree5),
    .dout108(r748tomtree5),
    .dout109(r749tomtree5),
    .dout110(r750tomtree5),
    .dout111(r751tomtree5),
    .dout112(r752tomtree5),
    .dout113(r753tomtree5),
    .dout114(r754tomtree5),
    .dout115(r755tomtree5),
    .dout116(r756tomtree5),
    .dout117(r757tomtree5),
    .dout118(r758tomtree5),
    .dout119(r759tomtree5),
    .dout120(r760tomtree5),
    .dout121(r761tomtree5),
    .dout122(r762tomtree5),
    .dout123(r763tomtree5),
    .dout124(r764tomtree5),
    .dout125(r765tomtree5),
    .dout126(r766tomtree5),
    .dout127(r767tomtree5)
  );

  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_6(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[6]),
    .din(mrgnsrcmuxout),
    .dout0(r768tomtree6),
    .dout1(r769tomtree6),
    .dout2(r770tomtree6),
    .dout3(r771tomtree6),
    .dout4(r772tomtree6),
    .dout5(r773tomtree6),
    .dout6(r774tomtree6),
    .dout7(r775tomtree6),
    .dout8(r776tomtree6),
    .dout9(r777tomtree6),
    .dout10(r778tomtree6),
    .dout11(r779tomtree6),
    .dout12(r780tomtree6),
    .dout13(r781tomtree6),
    .dout14(r782tomtree6),
    .dout15(r783tomtree6),
    .dout16(r784tomtree6),
    .dout17(r785tomtree6),
    .dout18(r786tomtree6),
    .dout19(r787tomtree6),
    .dout20(r788tomtree6),
    .dout21(r789tomtree6),
    .dout22(r790tomtree6),
    .dout23(r791tomtree6),
    .dout24(r792tomtree6),
    .dout25(r793tomtree6),
    .dout26(r794tomtree6),
    .dout27(r795tomtree6),
    .dout28(r796tomtree6),
    .dout29(r797tomtree6),
    .dout30(r798tomtree6),
    .dout31(r799tomtree6),
    .dout32(r800tomtree6),
    .dout33(r801tomtree6),
    .dout34(r802tomtree6),
    .dout35(r803tomtree6),
    .dout36(r804tomtree6),
    .dout37(r805tomtree6),
    .dout38(r806tomtree6),
    .dout39(r807tomtree6),
    .dout40(r808tomtree6),
    .dout41(r809tomtree6),
    .dout42(r810tomtree6),
    .dout43(r811tomtree6),
    .dout44(r812tomtree6),
    .dout45(r813tomtree6),
    .dout46(r814tomtree6),
    .dout47(r815tomtree6),
    .dout48(r816tomtree6),
    .dout49(r817tomtree6),
    .dout50(r818tomtree6),
    .dout51(r819tomtree6),
    .dout52(r820tomtree6),
    .dout53(r821tomtree6),
    .dout54(r822tomtree6),
    .dout55(r823tomtree6),
    .dout56(r824tomtree6),
    .dout57(r825tomtree6),
    .dout58(r826tomtree6),
    .dout59(r827tomtree6),
    .dout60(r828tomtree6),
    .dout61(r829tomtree6),
    .dout62(r830tomtree6),
    .dout63(r831tomtree6),
    .dout64(r832tomtree6),
    .dout65(r833tomtree6),
    .dout66(r834tomtree6),
    .dout67(r835tomtree6),
    .dout68(r836tomtree6),
    .dout69(r837tomtree6),
    .dout70(r838tomtree6),
    .dout71(r839tomtree6),
    .dout72(r840tomtree6),
    .dout73(r841tomtree6),
    .dout74(r842tomtree6),
    .dout75(r843tomtree6),
    .dout76(r844tomtree6),
    .dout77(r845tomtree6),
    .dout78(r846tomtree6),
    .dout79(r847tomtree6),
    .dout80(r848tomtree6),
    .dout81(r849tomtree6),
    .dout82(r850tomtree6),
    .dout83(r851tomtree6),
    .dout84(r852tomtree6),
    .dout85(r853tomtree6),
    .dout86(r854tomtree6),
    .dout87(r855tomtree6),
    .dout88(r856tomtree6),
    .dout89(r857tomtree6),
    .dout90(r858tomtree6),
    .dout91(r859tomtree6),
    .dout92(r860tomtree6),
    .dout93(r861tomtree6),
    .dout94(r862tomtree6),
    .dout95(r863tomtree6),
    .dout96(r864tomtree6),
    .dout97(r865tomtree6),
    .dout98(r866tomtree6),
    .dout99(r867tomtree6),
    .dout100(r868tomtree6),
    .dout101(r869tomtree6),
    .dout102(r870tomtree6),
    .dout103(r871tomtree6),
    .dout104(r872tomtree6),
    .dout105(r873tomtree6),
    .dout106(r874tomtree6),
    .dout107(r875tomtree6),
    .dout108(r876tomtree6),
    .dout109(r877tomtree6),
    .dout110(r878tomtree6),
    .dout111(r879tomtree6),
    .dout112(r880tomtree6),
    .dout113(r881tomtree6),
    .dout114(r882tomtree6),
    .dout115(r883tomtree6),
    .dout116(r884tomtree6),
    .dout117(r885tomtree6),
    .dout118(r886tomtree6),
    .dout119(r887tomtree6),
    .dout120(r888tomtree6),
    .dout121(r889tomtree6),
    .dout122(r890tomtree6),
    .dout123(r891tomtree6),
    .dout124(r892tomtree6),
    .dout125(r893tomtree6),
    .dout126(r894tomtree6),
    .dout127(r895tomtree6)
  );

  registers128 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_7(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[7]),
    .din(mrgnsrcmuxout),
    .dout0(r896tomtree7),
    .dout1(r897tomtree7),
    .dout2(r898tomtree7),
    .dout3(r899tomtree7),
    .dout4(r900tomtree7),
    .dout5(r901tomtree7),
    .dout6(r902tomtree7),
    .dout7(r903tomtree7),
    .dout8(r904tomtree7),
    .dout9(r905tomtree7),
    .dout10(r906tomtree7),
    .dout11(r907tomtree7),
    .dout12(r908tomtree7),
    .dout13(r909tomtree7),
    .dout14(r910tomtree7),
    .dout15(r911tomtree7),
    .dout16(r912tomtree7),
    .dout17(r913tomtree7),
    .dout18(r914tomtree7),
    .dout19(r915tomtree7),
    .dout20(r916tomtree7),
    .dout21(r917tomtree7),
    .dout22(r918tomtree7),
    .dout23(r919tomtree7),
    .dout24(r920tomtree7),
    .dout25(r921tomtree7),
    .dout26(r922tomtree7),
    .dout27(r923tomtree7),
    .dout28(r924tomtree7),
    .dout29(r925tomtree7),
    .dout30(r926tomtree7),
    .dout31(r927tomtree7),
    .dout32(r928tomtree7),
    .dout33(r929tomtree7),
    .dout34(r930tomtree7),
    .dout35(r931tomtree7),
    .dout36(r932tomtree7),
    .dout37(r933tomtree7),
    .dout38(r934tomtree7),
    .dout39(r935tomtree7),
    .dout40(r936tomtree7),
    .dout41(r937tomtree7),
    .dout42(r938tomtree7),
    .dout43(r939tomtree7),
    .dout44(r940tomtree7),
    .dout45(r941tomtree7),
    .dout46(r942tomtree7),
    .dout47(r943tomtree7),
    .dout48(r944tomtree7),
    .dout49(r945tomtree7),
    .dout50(r946tomtree7),
    .dout51(r947tomtree7),
    .dout52(r948tomtree7),
    .dout53(r949tomtree7),
    .dout54(r950tomtree7),
    .dout55(r951tomtree7),
    .dout56(r952tomtree7),
    .dout57(r953tomtree7),
    .dout58(r954tomtree7),
    .dout59(r955tomtree7),
    .dout60(r956tomtree7),
    .dout61(r957tomtree7),
    .dout62(r958tomtree7),
    .dout63(r959tomtree7),
    .dout64(r960tomtree7),
    .dout65(r961tomtree7),
    .dout66(r962tomtree7),
    .dout67(r963tomtree7),
    .dout68(r964tomtree7),
    .dout69(r965tomtree7),
    .dout70(r966tomtree7),
    .dout71(r967tomtree7),
    .dout72(r968tomtree7),
    .dout73(r969tomtree7),
    .dout74(r970tomtree7),
    .dout75(r971tomtree7),
    .dout76(r972tomtree7),
    .dout77(r973tomtree7),
    .dout78(r974tomtree7),
    .dout79(r975tomtree7),
    .dout80(r976tomtree7),
    .dout81(r977tomtree7),
    .dout82(r978tomtree7),
    .dout83(r979tomtree7),
    .dout84(r980tomtree7),
    .dout85(r981tomtree7),
    .dout86(r982tomtree7),
    .dout87(r983tomtree7),
    .dout88(r984tomtree7),
    .dout89(r985tomtree7),
    .dout90(r986tomtree7),
    .dout91(r987tomtree7),
    .dout92(r988tomtree7),
    .dout93(r989tomtree7),
    .dout94(r990tomtree7),
    .dout95(r991tomtree7),
    .dout96(r992tomtree7),
    .dout97(r993tomtree7),
    .dout98(r994tomtree7),
    .dout99(r995tomtree7),
    .dout100(r996tomtree7),
    .dout101(r997tomtree7),
    .dout102(r998tomtree7),
    .dout103(r999tomtree7),
    .dout104(r1000tomtree7),
    .dout105(r1001tomtree7),
    .dout106(r1002tomtree7),
    .dout107(r1003tomtree7),
    .dout108(r1004tomtree7),
    .dout109(r1005tomtree7),
    .dout110(r1006tomtree7),
    .dout111(r1007tomtree7),
    .dout112(r1008tomtree7),
    .dout113(r1009tomtree7),
    .dout114(r1010tomtree7),
    .dout115(r1011tomtree7),
    .dout116(r1012tomtree7),
    .dout117(r1013tomtree7),
    .dout118(r1014tomtree7),
    .dout119(r1015tomtree7),
    .dout120(r1016tomtree7),
    .dout121(r1017tomtree7),
    .dout122(r1018tomtree7),
    .dout123(r1019tomtree7),
    .dout124(r1020tomtree7),
    .dout125(r1021tomtree7),
    .dout126(r1022tomtree7),
    .dout127(r1023tomtree7)
  );
  
  mux2 #(.DATA_WIDTH(N_REGISTERSBANKS)) TrigMTreeSrcMux(
    .din0('b0), 
    .din1(decrb), 
    .sel(trigmtree), 
    .dout(trigmtreesrcmuxout)
  );
  
  register #(.DATA_WIDTH(N_REGISTERSBANKS)) RTrigMTreeSrcMux(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(trigmtreesrcmuxout),
    .dout(trigmtreeold)
  );
  
  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_0(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[0]),
    .din0(r0tomtree0),
    .din1(r1tomtree0),
    .din2(r2tomtree0),
    .din3(r3tomtree0),
    .din4(r4tomtree0),
    .din5(r5tomtree0),
    .din6(r6tomtree0),
    .din7(r7tomtree0),
    .din8(r8tomtree0),
    .din9(r9tomtree0),
    .din10(r10tomtree0),
    .din11(r11tomtree0),
    .din12(r12tomtree0),
    .din13(r13tomtree0),
    .din14(r14tomtree0),
    .din15(r15tomtree0),
    .din16(r16tomtree0),
    .din17(r17tomtree0),
    .din18(r18tomtree0),
    .din19(r19tomtree0),
    .din20(r20tomtree0),
    .din21(r21tomtree0),
    .din22(r22tomtree0),
    .din23(r23tomtree0),
    .din24(r24tomtree0),
    .din25(r25tomtree0),
    .din26(r26tomtree0),
    .din27(r27tomtree0),
    .din28(r28tomtree0),
    .din29(r29tomtree0),
    .din30(r30tomtree0),
    .din31(r31tomtree0),
    .din32(r32tomtree0),
    .din33(r33tomtree0),
    .din34(r34tomtree0),
    .din35(r35tomtree0),
    .din36(r36tomtree0),
    .din37(r37tomtree0),
    .din38(r38tomtree0),
    .din39(r39tomtree0),
    .din40(r40tomtree0),
    .din41(r41tomtree0),
    .din42(r42tomtree0),
    .din43(r43tomtree0),
    .din44(r44tomtree0),
    .din45(r45tomtree0),
    .din46(r46tomtree0),
    .din47(r47tomtree0),
    .din48(r48tomtree0),
    .din49(r49tomtree0),
    .din50(r50tomtree0),
    .din51(r51tomtree0),
    .din52(r52tomtree0),
    .din53(r53tomtree0),
    .din54(r54tomtree0),
    .din55(r55tomtree0),
    .din56(r56tomtree0),
    .din57(r57tomtree0),
    .din58(r58tomtree0),
    .din59(r59tomtree0),
    .din60(r60tomtree0),
    .din61(r61tomtree0),
    .din62(r62tomtree0),
    .din63(r63tomtree0),
    .din64(r64tomtree0),
    .din65(r65tomtree0),
    .din66(r66tomtree0),
    .din67(r67tomtree0),
    .din68(r68tomtree0),
    .din69(r69tomtree0),
    .din70(r70tomtree0),
    .din71(r71tomtree0),
    .din72(r72tomtree0),
    .din73(r73tomtree0),
    .din74(r74tomtree0),
    .din75(r75tomtree0),
    .din76(r76tomtree0),
    .din77(r77tomtree0),
    .din78(r78tomtree0),
    .din79(r79tomtree0),
    .din80(r80tomtree0),
    .din81(r81tomtree0),
    .din82(r82tomtree0),
    .din83(r83tomtree0),
    .din84(r84tomtree0),
    .din85(r85tomtree0),
    .din86(r86tomtree0),
    .din87(r87tomtree0),
    .din88(r88tomtree0),
    .din89(r89tomtree0),
    .din90(r90tomtree0),
    .din91(r91tomtree0),
    .din92(r92tomtree0),
    .din93(r93tomtree0),
    .din94(r94tomtree0),
    .din95(r95tomtree0),
    .din96(r96tomtree0),
    .din97(r97tomtree0),
    .din98(r98tomtree0),
    .din99(r99tomtree0),
    .din100(r100tomtree0),
    .din101(r101tomtree0),
    .din102(r102tomtree0),
    .din103(r103tomtree0),
    .din104(r104tomtree0),
    .din105(r105tomtree0),
    .din106(r106tomtree0),
    .din107(r107tomtree0),
    .din108(r108tomtree0),
    .din109(r109tomtree0),
    .din110(r110tomtree0),
    .din111(r111tomtree0),
    .din112(r112tomtree0),
    .din113(r113tomtree0),
    .din114(r114tomtree0),
    .din115(r115tomtree0),
    .din116(r116tomtree0),
    .din117(r117tomtree0),
    .din118(r118tomtree0),
    .din119(r119tomtree0),
    .din120(r120tomtree0),
    .din121(r121tomtree0),
    .din122(r122tomtree0),
    .din123(r123tomtree0),
    .din124(r124tomtree0),
    .din125(r125tomtree0),
    .din126(r126tomtree0),
    .din127(r127tomtree0),
    .max(mtree0tomaxsrcmux)
  );

  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_1(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[1]),
    .din0(r128tomtree1),
    .din1(r129tomtree1),
    .din2(r130tomtree1),
    .din3(r131tomtree1),
    .din4(r132tomtree1),
    .din5(r133tomtree1),
    .din6(r134tomtree1),
    .din7(r135tomtree1),
    .din8(r136tomtree1),
    .din9(r137tomtree1),
    .din10(r138tomtree1),
    .din11(r139tomtree1),
    .din12(r140tomtree1),
    .din13(r141tomtree1),
    .din14(r142tomtree1),
    .din15(r143tomtree1),
    .din16(r144tomtree1),
    .din17(r145tomtree1),
    .din18(r146tomtree1),
    .din19(r147tomtree1),
    .din20(r148tomtree1),
    .din21(r149tomtree1),
    .din22(r150tomtree1),
    .din23(r151tomtree1),
    .din24(r152tomtree1),
    .din25(r153tomtree1),
    .din26(r154tomtree1),
    .din27(r155tomtree1),
    .din28(r156tomtree1),
    .din29(r157tomtree1),
    .din30(r158tomtree1),
    .din31(r159tomtree1),
    .din32(r160tomtree1),
    .din33(r161tomtree1),
    .din34(r162tomtree1),
    .din35(r163tomtree1),
    .din36(r164tomtree1),
    .din37(r165tomtree1),
    .din38(r166tomtree1),
    .din39(r167tomtree1),
    .din40(r168tomtree1),
    .din41(r169tomtree1),
    .din42(r170tomtree1),
    .din43(r171tomtree1),
    .din44(r172tomtree1),
    .din45(r173tomtree1),
    .din46(r174tomtree1),
    .din47(r175tomtree1),
    .din48(r176tomtree1),
    .din49(r177tomtree1),
    .din50(r178tomtree1),
    .din51(r179tomtree1),
    .din52(r180tomtree1),
    .din53(r181tomtree1),
    .din54(r182tomtree1),
    .din55(r183tomtree1),
    .din56(r184tomtree1),
    .din57(r185tomtree1),
    .din58(r186tomtree1),
    .din59(r187tomtree1),
    .din60(r188tomtree1),
    .din61(r189tomtree1),
    .din62(r190tomtree1),
    .din63(r191tomtree1),
    .din64(r192tomtree1),
    .din65(r193tomtree1),
    .din66(r194tomtree1),
    .din67(r195tomtree1),
    .din68(r196tomtree1),
    .din69(r197tomtree1),
    .din70(r198tomtree1),
    .din71(r199tomtree1),
    .din72(r200tomtree1),
    .din73(r201tomtree1),
    .din74(r202tomtree1),
    .din75(r203tomtree1),
    .din76(r204tomtree1),
    .din77(r205tomtree1),
    .din78(r206tomtree1),
    .din79(r207tomtree1),
    .din80(r208tomtree1),
    .din81(r209tomtree1),
    .din82(r210tomtree1),
    .din83(r211tomtree1),
    .din84(r212tomtree1),
    .din85(r213tomtree1),
    .din86(r214tomtree1),
    .din87(r215tomtree1),
    .din88(r216tomtree1),
    .din89(r217tomtree1),
    .din90(r218tomtree1),
    .din91(r219tomtree1),
    .din92(r220tomtree1),
    .din93(r221tomtree1),
    .din94(r222tomtree1),
    .din95(r223tomtree1),
    .din96(r224tomtree1),
    .din97(r225tomtree1),
    .din98(r226tomtree1),
    .din99(r227tomtree1),
    .din100(r228tomtree1),
    .din101(r229tomtree1),
    .din102(r230tomtree1),
    .din103(r231tomtree1),
    .din104(r232tomtree1),
    .din105(r233tomtree1),
    .din106(r234tomtree1),
    .din107(r235tomtree1),
    .din108(r236tomtree1),
    .din109(r237tomtree1),
    .din110(r238tomtree1),
    .din111(r239tomtree1),
    .din112(r240tomtree1),
    .din113(r241tomtree1),
    .din114(r242tomtree1),
    .din115(r243tomtree1),
    .din116(r244tomtree1),
    .din117(r245tomtree1),
    .din118(r246tomtree1),
    .din119(r247tomtree1),
    .din120(r248tomtree1),
    .din121(r249tomtree1),
    .din122(r250tomtree1),
    .din123(r251tomtree1),
    .din124(r252tomtree1),
    .din125(r253tomtree1),
    .din126(r254tomtree1),
    .din127(r255tomtree1),
    .max(mtree1tomaxsrcmux)
  );

  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_2(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[2]),
    .din0(r256tomtree2),
    .din1(r257tomtree2),
    .din2(r258tomtree2),
    .din3(r259tomtree2),
    .din4(r260tomtree2),
    .din5(r261tomtree2),
    .din6(r262tomtree2),
    .din7(r263tomtree2),
    .din8(r264tomtree2),
    .din9(r265tomtree2),
    .din10(r266tomtree2),
    .din11(r267tomtree2),
    .din12(r268tomtree2),
    .din13(r269tomtree2),
    .din14(r270tomtree2),
    .din15(r271tomtree2),
    .din16(r272tomtree2),
    .din17(r273tomtree2),
    .din18(r274tomtree2),
    .din19(r275tomtree2),
    .din20(r276tomtree2),
    .din21(r277tomtree2),
    .din22(r278tomtree2),
    .din23(r279tomtree2),
    .din24(r280tomtree2),
    .din25(r281tomtree2),
    .din26(r282tomtree2),
    .din27(r283tomtree2),
    .din28(r284tomtree2),
    .din29(r285tomtree2),
    .din30(r286tomtree2),
    .din31(r287tomtree2),
    .din32(r288tomtree2),
    .din33(r289tomtree2),
    .din34(r290tomtree2),
    .din35(r291tomtree2),
    .din36(r292tomtree2),
    .din37(r293tomtree2),
    .din38(r294tomtree2),
    .din39(r295tomtree2),
    .din40(r296tomtree2),
    .din41(r297tomtree2),
    .din42(r298tomtree2),
    .din43(r299tomtree2),
    .din44(r300tomtree2),
    .din45(r301tomtree2),
    .din46(r302tomtree2),
    .din47(r303tomtree2),
    .din48(r304tomtree2),
    .din49(r305tomtree2),
    .din50(r306tomtree2),
    .din51(r307tomtree2),
    .din52(r308tomtree2),
    .din53(r309tomtree2),
    .din54(r310tomtree2),
    .din55(r311tomtree2),
    .din56(r312tomtree2),
    .din57(r313tomtree2),
    .din58(r314tomtree2),
    .din59(r315tomtree2),
    .din60(r316tomtree2),
    .din61(r317tomtree2),
    .din62(r318tomtree2),
    .din63(r319tomtree2),
    .din64(r320tomtree2),
    .din65(r321tomtree2),
    .din66(r322tomtree2),
    .din67(r323tomtree2),
    .din68(r324tomtree2),
    .din69(r325tomtree2),
    .din70(r326tomtree2),
    .din71(r327tomtree2),
    .din72(r328tomtree2),
    .din73(r329tomtree2),
    .din74(r330tomtree2),
    .din75(r331tomtree2),
    .din76(r332tomtree2),
    .din77(r333tomtree2),
    .din78(r334tomtree2),
    .din79(r335tomtree2),
    .din80(r336tomtree2),
    .din81(r337tomtree2),
    .din82(r338tomtree2),
    .din83(r339tomtree2),
    .din84(r340tomtree2),
    .din85(r341tomtree2),
    .din86(r342tomtree2),
    .din87(r343tomtree2),
    .din88(r344tomtree2),
    .din89(r345tomtree2),
    .din90(r346tomtree2),
    .din91(r347tomtree2),
    .din92(r348tomtree2),
    .din93(r349tomtree2),
    .din94(r350tomtree2),
    .din95(r351tomtree2),
    .din96(r352tomtree2),
    .din97(r353tomtree2),
    .din98(r354tomtree2),
    .din99(r355tomtree2),
    .din100(r356tomtree2),
    .din101(r357tomtree2),
    .din102(r358tomtree2),
    .din103(r359tomtree2),
    .din104(r360tomtree2),
    .din105(r361tomtree2),
    .din106(r362tomtree2),
    .din107(r363tomtree2),
    .din108(r364tomtree2),
    .din109(r365tomtree2),
    .din110(r366tomtree2),
    .din111(r367tomtree2),
    .din112(r368tomtree2),
    .din113(r369tomtree2),
    .din114(r370tomtree2),
    .din115(r371tomtree2),
    .din116(r372tomtree2),
    .din117(r373tomtree2),
    .din118(r374tomtree2),
    .din119(r375tomtree2),
    .din120(r376tomtree2),
    .din121(r377tomtree2),
    .din122(r378tomtree2),
    .din123(r379tomtree2),
    .din124(r380tomtree2),
    .din125(r381tomtree2),
    .din126(r382tomtree2),
    .din127(r383tomtree2),
    .max(mtree2tomaxsrcmux)
  );

  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_3(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[3]),
    .din0(r384tomtree3),
    .din1(r385tomtree3),
    .din2(r386tomtree3),
    .din3(r387tomtree3),
    .din4(r388tomtree3),
    .din5(r389tomtree3),
    .din6(r390tomtree3),
    .din7(r391tomtree3),
    .din8(r392tomtree3),
    .din9(r393tomtree3),
    .din10(r394tomtree3),
    .din11(r395tomtree3),
    .din12(r396tomtree3),
    .din13(r397tomtree3),
    .din14(r398tomtree3),
    .din15(r399tomtree3),
    .din16(r400tomtree3),
    .din17(r401tomtree3),
    .din18(r402tomtree3),
    .din19(r403tomtree3),
    .din20(r404tomtree3),
    .din21(r405tomtree3),
    .din22(r406tomtree3),
    .din23(r407tomtree3),
    .din24(r408tomtree3),
    .din25(r409tomtree3),
    .din26(r410tomtree3),
    .din27(r411tomtree3),
    .din28(r412tomtree3),
    .din29(r413tomtree3),
    .din30(r414tomtree3),
    .din31(r415tomtree3),
    .din32(r416tomtree3),
    .din33(r417tomtree3),
    .din34(r418tomtree3),
    .din35(r419tomtree3),
    .din36(r420tomtree3),
    .din37(r421tomtree3),
    .din38(r422tomtree3),
    .din39(r423tomtree3),
    .din40(r424tomtree3),
    .din41(r425tomtree3),
    .din42(r426tomtree3),
    .din43(r427tomtree3),
    .din44(r428tomtree3),
    .din45(r429tomtree3),
    .din46(r430tomtree3),
    .din47(r431tomtree3),
    .din48(r432tomtree3),
    .din49(r433tomtree3),
    .din50(r434tomtree3),
    .din51(r435tomtree3),
    .din52(r436tomtree3),
    .din53(r437tomtree3),
    .din54(r438tomtree3),
    .din55(r439tomtree3),
    .din56(r440tomtree3),
    .din57(r441tomtree3),
    .din58(r442tomtree3),
    .din59(r443tomtree3),
    .din60(r444tomtree3),
    .din61(r445tomtree3),
    .din62(r446tomtree3),
    .din63(r447tomtree3),
    .din64(r448tomtree3),
    .din65(r449tomtree3),
    .din66(r450tomtree3),
    .din67(r451tomtree3),
    .din68(r452tomtree3),
    .din69(r453tomtree3),
    .din70(r454tomtree3),
    .din71(r455tomtree3),
    .din72(r456tomtree3),
    .din73(r457tomtree3),
    .din74(r458tomtree3),
    .din75(r459tomtree3),
    .din76(r460tomtree3),
    .din77(r461tomtree3),
    .din78(r462tomtree3),
    .din79(r463tomtree3),
    .din80(r464tomtree3),
    .din81(r465tomtree3),
    .din82(r466tomtree3),
    .din83(r467tomtree3),
    .din84(r468tomtree3),
    .din85(r469tomtree3),
    .din86(r470tomtree3),
    .din87(r471tomtree3),
    .din88(r472tomtree3),
    .din89(r473tomtree3),
    .din90(r474tomtree3),
    .din91(r475tomtree3),
    .din92(r476tomtree3),
    .din93(r477tomtree3),
    .din94(r478tomtree3),
    .din95(r479tomtree3),
    .din96(r480tomtree3),
    .din97(r481tomtree3),
    .din98(r482tomtree3),
    .din99(r483tomtree3),
    .din100(r484tomtree3),
    .din101(r485tomtree3),
    .din102(r486tomtree3),
    .din103(r487tomtree3),
    .din104(r488tomtree3),
    .din105(r489tomtree3),
    .din106(r490tomtree3),
    .din107(r491tomtree3),
    .din108(r492tomtree3),
    .din109(r493tomtree3),
    .din110(r494tomtree3),
    .din111(r495tomtree3),
    .din112(r496tomtree3),
    .din113(r497tomtree3),
    .din114(r498tomtree3),
    .din115(r499tomtree3),
    .din116(r500tomtree3),
    .din117(r501tomtree3),
    .din118(r502tomtree3),
    .din119(r503tomtree3),
    .din120(r504tomtree3),
    .din121(r505tomtree3),
    .din122(r506tomtree3),
    .din123(r507tomtree3),
    .din124(r508tomtree3),
    .din125(r509tomtree3),
    .din126(r510tomtree3),
    .din127(r511tomtree3),
    .max(mtree3tomaxsrcmux)
  );
  
  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_4(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[4]),
    .din0(r512tomtree4),
    .din1(r513tomtree4),
    .din2(r514tomtree4),
    .din3(r515tomtree4),
    .din4(r516tomtree4),
    .din5(r517tomtree4),
    .din6(r518tomtree4),
    .din7(r519tomtree4),
    .din8(r520tomtree4),
    .din9(r521tomtree4),
    .din10(r522tomtree4),
    .din11(r523tomtree4),
    .din12(r524tomtree4),
    .din13(r525tomtree4),
    .din14(r526tomtree4),
    .din15(r527tomtree4),
    .din16(r528tomtree4),
    .din17(r529tomtree4),
    .din18(r530tomtree4),
    .din19(r531tomtree4),
    .din20(r532tomtree4),
    .din21(r533tomtree4),
    .din22(r534tomtree4),
    .din23(r535tomtree4),
    .din24(r536tomtree4),
    .din25(r537tomtree4),
    .din26(r538tomtree4),
    .din27(r539tomtree4),
    .din28(r540tomtree4),
    .din29(r541tomtree4),
    .din30(r542tomtree4),
    .din31(r543tomtree4),
    .din32(r544tomtree4),
    .din33(r545tomtree4),
    .din34(r546tomtree4),
    .din35(r547tomtree4),
    .din36(r548tomtree4),
    .din37(r549tomtree4),
    .din38(r550tomtree4),
    .din39(r551tomtree4),
    .din40(r552tomtree4),
    .din41(r553tomtree4),
    .din42(r554tomtree4),
    .din43(r555tomtree4),
    .din44(r556tomtree4),
    .din45(r557tomtree4),
    .din46(r558tomtree4),
    .din47(r559tomtree4),
    .din48(r560tomtree4),
    .din49(r561tomtree4),
    .din50(r562tomtree4),
    .din51(r563tomtree4),
    .din52(r564tomtree4),
    .din53(r565tomtree4),
    .din54(r566tomtree4),
    .din55(r567tomtree4),
    .din56(r568tomtree4),
    .din57(r569tomtree4),
    .din58(r570tomtree4),
    .din59(r571tomtree4),
    .din60(r572tomtree4),
    .din61(r573tomtree4),
    .din62(r574tomtree4),
    .din63(r575tomtree4),
    .din64(r576tomtree4),
    .din65(r577tomtree4),
    .din66(r578tomtree4),
    .din67(r579tomtree4),
    .din68(r580tomtree4),
    .din69(r581tomtree4),
    .din70(r582tomtree4),
    .din71(r583tomtree4),
    .din72(r584tomtree4),
    .din73(r585tomtree4),
    .din74(r586tomtree4),
    .din75(r587tomtree4),
    .din76(r588tomtree4),
    .din77(r589tomtree4),
    .din78(r590tomtree4),
    .din79(r591tomtree4),
    .din80(r592tomtree4),
    .din81(r593tomtree4),
    .din82(r594tomtree4),
    .din83(r595tomtree4),
    .din84(r596tomtree4),
    .din85(r597tomtree4),
    .din86(r598tomtree4),
    .din87(r599tomtree4),
    .din88(r600tomtree4),
    .din89(r601tomtree4),
    .din90(r602tomtree4),
    .din91(r603tomtree4),
    .din92(r604tomtree4),
    .din93(r605tomtree4),
    .din94(r606tomtree4),
    .din95(r607tomtree4),
    .din96(r608tomtree4),
    .din97(r609tomtree4),
    .din98(r610tomtree4),
    .din99(r611tomtree4),
    .din100(r612tomtree4),
    .din101(r613tomtree4),
    .din102(r614tomtree4),
    .din103(r615tomtree4),
    .din104(r616tomtree4),
    .din105(r617tomtree4),
    .din106(r618tomtree4),
    .din107(r619tomtree4),
    .din108(r620tomtree4),
    .din109(r621tomtree4),
    .din110(r622tomtree4),
    .din111(r623tomtree4),
    .din112(r624tomtree4),
    .din113(r625tomtree4),
    .din114(r626tomtree4),
    .din115(r627tomtree4),
    .din116(r628tomtree4),
    .din117(r629tomtree4),
    .din118(r630tomtree4),
    .din119(r631tomtree4),
    .din120(r632tomtree4),
    .din121(r633tomtree4),
    .din122(r634tomtree4),
    .din123(r635tomtree4),
    .din124(r636tomtree4),
    .din125(r637tomtree4),
    .din126(r638tomtree4),
    .din127(r639tomtree4),
    .max(mtree4tomaxsrcmux)
  );

  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_5(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[5]),
    .din0(r640tomtree5),
    .din1(r641tomtree5),
    .din2(r642tomtree5),
    .din3(r643tomtree5),
    .din4(r644tomtree5),
    .din5(r645tomtree5),
    .din6(r646tomtree5),
    .din7(r647tomtree5),
    .din8(r648tomtree5),
    .din9(r649tomtree5),
    .din10(r650tomtree5),
    .din11(r651tomtree5),
    .din12(r652tomtree5),
    .din13(r653tomtree5),
    .din14(r654tomtree5),
    .din15(r655tomtree5),
    .din16(r656tomtree5),
    .din17(r657tomtree5),
    .din18(r658tomtree5),
    .din19(r659tomtree5),
    .din20(r660tomtree5),
    .din21(r661tomtree5),
    .din22(r662tomtree5),
    .din23(r663tomtree5),
    .din24(r664tomtree5),
    .din25(r665tomtree5),
    .din26(r666tomtree5),
    .din27(r667tomtree5),
    .din28(r668tomtree5),
    .din29(r669tomtree5),
    .din30(r670tomtree5),
    .din31(r671tomtree5),
    .din32(r672tomtree5),
    .din33(r673tomtree5),
    .din34(r674tomtree5),
    .din35(r675tomtree5),
    .din36(r676tomtree5),
    .din37(r677tomtree5),
    .din38(r678tomtree5),
    .din39(r679tomtree5),
    .din40(r680tomtree5),
    .din41(r681tomtree5),
    .din42(r682tomtree5),
    .din43(r683tomtree5),
    .din44(r684tomtree5),
    .din45(r685tomtree5),
    .din46(r686tomtree5),
    .din47(r687tomtree5),
    .din48(r688tomtree5),
    .din49(r689tomtree5),
    .din50(r690tomtree5),
    .din51(r691tomtree5),
    .din52(r692tomtree5),
    .din53(r693tomtree5),
    .din54(r694tomtree5),
    .din55(r695tomtree5),
    .din56(r696tomtree5),
    .din57(r697tomtree5),
    .din58(r698tomtree5),
    .din59(r699tomtree5),
    .din60(r700tomtree5),
    .din61(r701tomtree5),
    .din62(r702tomtree5),
    .din63(r703tomtree5),
    .din64(r704tomtree5),
    .din65(r705tomtree5),
    .din66(r706tomtree5),
    .din67(r707tomtree5),
    .din68(r708tomtree5),
    .din69(r709tomtree5),
    .din70(r710tomtree5),
    .din71(r711tomtree5),
    .din72(r712tomtree5),
    .din73(r713tomtree5),
    .din74(r714tomtree5),
    .din75(r715tomtree5),
    .din76(r716tomtree5),
    .din77(r717tomtree5),
    .din78(r718tomtree5),
    .din79(r719tomtree5),
    .din80(r720tomtree5),
    .din81(r721tomtree5),
    .din82(r722tomtree5),
    .din83(r723tomtree5),
    .din84(r724tomtree5),
    .din85(r725tomtree5),
    .din86(r726tomtree5),
    .din87(r727tomtree5),
    .din88(r728tomtree5),
    .din89(r729tomtree5),
    .din90(r730tomtree5),
    .din91(r731tomtree5),
    .din92(r732tomtree5),
    .din93(r733tomtree5),
    .din94(r734tomtree5),
    .din95(r735tomtree5),
    .din96(r736tomtree5),
    .din97(r737tomtree5),
    .din98(r738tomtree5),
    .din99(r739tomtree5),
    .din100(r740tomtree5),
    .din101(r741tomtree5),
    .din102(r742tomtree5),
    .din103(r743tomtree5),
    .din104(r744tomtree5),
    .din105(r745tomtree5),
    .din106(r746tomtree5),
    .din107(r747tomtree5),
    .din108(r748tomtree5),
    .din109(r749tomtree5),
    .din110(r750tomtree5),
    .din111(r751tomtree5),
    .din112(r752tomtree5),
    .din113(r753tomtree5),
    .din114(r754tomtree5),
    .din115(r755tomtree5),
    .din116(r756tomtree5),
    .din117(r757tomtree5),
    .din118(r758tomtree5),
    .din119(r759tomtree5),
    .din120(r760tomtree5),
    .din121(r761tomtree5),
    .din122(r762tomtree5),
    .din123(r763tomtree5),
    .din124(r764tomtree5),
    .din125(r765tomtree5),
    .din126(r766tomtree5),
    .din127(r767tomtree5),
    .max(mtree5tomaxsrcmux)
  );

  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_6(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[6]),
    .din0(r768tomtree6),
    .din1(r769tomtree6),
    .din2(r770tomtree6),
    .din3(r771tomtree6),
    .din4(r772tomtree6),
    .din5(r773tomtree6),
    .din6(r774tomtree6),
    .din7(r775tomtree6),
    .din8(r776tomtree6),
    .din9(r777tomtree6),
    .din10(r778tomtree6),
    .din11(r779tomtree6),
    .din12(r780tomtree6),
    .din13(r781tomtree6),
    .din14(r782tomtree6),
    .din15(r783tomtree6),
    .din16(r784tomtree6),
    .din17(r785tomtree6),
    .din18(r786tomtree6),
    .din19(r787tomtree6),
    .din20(r788tomtree6),
    .din21(r789tomtree6),
    .din22(r790tomtree6),
    .din23(r791tomtree6),
    .din24(r792tomtree6),
    .din25(r793tomtree6),
    .din26(r794tomtree6),
    .din27(r795tomtree6),
    .din28(r796tomtree6),
    .din29(r797tomtree6),
    .din30(r798tomtree6),
    .din31(r799tomtree6),
    .din32(r800tomtree6),
    .din33(r801tomtree6),
    .din34(r802tomtree6),
    .din35(r803tomtree6),
    .din36(r804tomtree6),
    .din37(r805tomtree6),
    .din38(r806tomtree6),
    .din39(r807tomtree6),
    .din40(r808tomtree6),
    .din41(r809tomtree6),
    .din42(r810tomtree6),
    .din43(r811tomtree6),
    .din44(r812tomtree6),
    .din45(r813tomtree6),
    .din46(r814tomtree6),
    .din47(r815tomtree6),
    .din48(r816tomtree6),
    .din49(r817tomtree6),
    .din50(r818tomtree6),
    .din51(r819tomtree6),
    .din52(r820tomtree6),
    .din53(r821tomtree6),
    .din54(r822tomtree6),
    .din55(r823tomtree6),
    .din56(r824tomtree6),
    .din57(r825tomtree6),
    .din58(r826tomtree6),
    .din59(r827tomtree6),
    .din60(r828tomtree6),
    .din61(r829tomtree6),
    .din62(r830tomtree6),
    .din63(r831tomtree6),
    .din64(r832tomtree6),
    .din65(r833tomtree6),
    .din66(r834tomtree6),
    .din67(r835tomtree6),
    .din68(r836tomtree6),
    .din69(r837tomtree6),
    .din70(r838tomtree6),
    .din71(r839tomtree6),
    .din72(r840tomtree6),
    .din73(r841tomtree6),
    .din74(r842tomtree6),
    .din75(r843tomtree6),
    .din76(r844tomtree6),
    .din77(r845tomtree6),
    .din78(r846tomtree6),
    .din79(r847tomtree6),
    .din80(r848tomtree6),
    .din81(r849tomtree6),
    .din82(r850tomtree6),
    .din83(r851tomtree6),
    .din84(r852tomtree6),
    .din85(r853tomtree6),
    .din86(r854tomtree6),
    .din87(r855tomtree6),
    .din88(r856tomtree6),
    .din89(r857tomtree6),
    .din90(r858tomtree6),
    .din91(r859tomtree6),
    .din92(r860tomtree6),
    .din93(r861tomtree6),
    .din94(r862tomtree6),
    .din95(r863tomtree6),
    .din96(r864tomtree6),
    .din97(r865tomtree6),
    .din98(r866tomtree6),
    .din99(r867tomtree6),
    .din100(r868tomtree6),
    .din101(r869tomtree6),
    .din102(r870tomtree6),
    .din103(r871tomtree6),
    .din104(r872tomtree6),
    .din105(r873tomtree6),
    .din106(r874tomtree6),
    .din107(r875tomtree6),
    .din108(r876tomtree6),
    .din109(r877tomtree6),
    .din110(r878tomtree6),
    .din111(r879tomtree6),
    .din112(r880tomtree6),
    .din113(r881tomtree6),
    .din114(r882tomtree6),
    .din115(r883tomtree6),
    .din116(r884tomtree6),
    .din117(r885tomtree6),
    .din118(r886tomtree6),
    .din119(r887tomtree6),
    .din120(r888tomtree6),
    .din121(r889tomtree6),
    .din122(r890tomtree6),
    .din123(r891tomtree6),
    .din124(r892tomtree6),
    .din125(r893tomtree6),
    .din126(r894tomtree6),
    .din127(r895tomtree6),
    .max(mtree6tomaxsrcmux)
  );

  maxtree128 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_7(
    .clk(clk),
    .rst_n(rst_n),
    .start(trigmtreeold[7]),
    .din0(r896tomtree7),
    .din1(r897tomtree7),
    .din2(r898tomtree7),
    .din3(r899tomtree7),
    .din4(r900tomtree7),
    .din5(r901tomtree7),
    .din6(r902tomtree7),
    .din7(r903tomtree7),
    .din8(r904tomtree7),
    .din9(r905tomtree7),
    .din10(r906tomtree7),
    .din11(r907tomtree7),
    .din12(r908tomtree7),
    .din13(r909tomtree7),
    .din14(r910tomtree7),
    .din15(r911tomtree7),
    .din16(r912tomtree7),
    .din17(r913tomtree7),
    .din18(r914tomtree7),
    .din19(r915tomtree7),
    .din20(r916tomtree7),
    .din21(r917tomtree7),
    .din22(r918tomtree7),
    .din23(r919tomtree7),
    .din24(r920tomtree7),
    .din25(r921tomtree7),
    .din26(r922tomtree7),
    .din27(r923tomtree7),
    .din28(r924tomtree7),
    .din29(r925tomtree7),
    .din30(r926tomtree7),
    .din31(r927tomtree7),
    .din32(r928tomtree7),
    .din33(r929tomtree7),
    .din34(r930tomtree7),
    .din35(r931tomtree7),
    .din36(r932tomtree7),
    .din37(r933tomtree7),
    .din38(r934tomtree7),
    .din39(r935tomtree7),
    .din40(r936tomtree7),
    .din41(r937tomtree7),
    .din42(r938tomtree7),
    .din43(r939tomtree7),
    .din44(r940tomtree7),
    .din45(r941tomtree7),
    .din46(r942tomtree7),
    .din47(r943tomtree7),
    .din48(r944tomtree7),
    .din49(r945tomtree7),
    .din50(r946tomtree7),
    .din51(r947tomtree7),
    .din52(r948tomtree7),
    .din53(r949tomtree7),
    .din54(r950tomtree7),
    .din55(r951tomtree7),
    .din56(r952tomtree7),
    .din57(r953tomtree7),
    .din58(r954tomtree7),
    .din59(r955tomtree7),
    .din60(r956tomtree7),
    .din61(r957tomtree7),
    .din62(r958tomtree7),
    .din63(r959tomtree7),
    .din64(r960tomtree7),
    .din65(r961tomtree7),
    .din66(r962tomtree7),
    .din67(r963tomtree7),
    .din68(r964tomtree7),
    .din69(r965tomtree7),
    .din70(r966tomtree7),
    .din71(r967tomtree7),
    .din72(r968tomtree7),
    .din73(r969tomtree7),
    .din74(r970tomtree7),
    .din75(r971tomtree7),
    .din76(r972tomtree7),
    .din77(r973tomtree7),
    .din78(r974tomtree7),
    .din79(r975tomtree7),
    .din80(r976tomtree7),
    .din81(r977tomtree7),
    .din82(r978tomtree7),
    .din83(r979tomtree7),
    .din84(r980tomtree7),
    .din85(r981tomtree7),
    .din86(r982tomtree7),
    .din87(r983tomtree7),
    .din88(r984tomtree7),
    .din89(r985tomtree7),
    .din90(r986tomtree7),
    .din91(r987tomtree7),
    .din92(r988tomtree7),
    .din93(r989tomtree7),
    .din94(r990tomtree7),
    .din95(r991tomtree7),
    .din96(r992tomtree7),
    .din97(r993tomtree7),
    .din98(r994tomtree7),
    .din99(r995tomtree7),
    .din100(r996tomtree7),
    .din101(r997tomtree7),
    .din102(r998tomtree7),
    .din103(r999tomtree7),
    .din104(r1000tomtree7),
    .din105(r1001tomtree7),
    .din106(r1002tomtree7),
    .din107(r1003tomtree7),
    .din108(r1004tomtree7),
    .din109(r1005tomtree7),
    .din110(r1006tomtree7),
    .din111(r1007tomtree7),
    .din112(r1008tomtree7),
    .din113(r1009tomtree7),
    .din114(r1010tomtree7),
    .din115(r1011tomtree7),
    .din116(r1012tomtree7),
    .din117(r1013tomtree7),
    .din118(r1014tomtree7),
    .din119(r1015tomtree7),
    .din120(r1016tomtree7),
    .din121(r1017tomtree7),
    .din122(r1018tomtree7),
    .din123(r1019tomtree7),
    .din124(r1020tomtree7),
    .din125(r1021tomtree7),
    .din126(r1022tomtree7),
    .din127(r1023tomtree7),
    .max(mtree7tomaxsrcmux)
  );
  
  mux8 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) MaxSrcMux(
    .din0(mtree0tomaxsrcmux),
    .din1(mtree1tomaxsrcmux),
    .din2(mtree2tomaxsrcmux),
    .din3(mtree3tomaxsrcmux),
    .din4(mtree4tomaxsrcmux),
    .din5(mtree5tomaxsrcmux),
    .din6(mtree6tomaxsrcmux),
    .din7(mtree7tomaxsrcmux),
    .sel(cntrb),
    .dout(maxsrcmuxtocmp)
  );

  comparator #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH), .N_REGISTERS(N_REGISTERS)) Cmp(
    .max(maxsrcmuxtocmp),
    .margin({mrgnindx,mrgn}),
    .trig(trigmax),
    .r_sel(rcmp),
    .dout(mrgncmp)
  );
  
  mux1024 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) OutSrcMux(
    .din0(r0tomtree0),
    .din1(r1tomtree0),
    .din2(r2tomtree0),
    .din3(r3tomtree0),
    .din4(r4tomtree0),
    .din5(r5tomtree0),
    .din6(r6tomtree0),
    .din7(r7tomtree0),
    .din8(r8tomtree0),
    .din9(r9tomtree0),
    .din10(r10tomtree0),
    .din11(r11tomtree0),
    .din12(r12tomtree0),
    .din13(r13tomtree0),
    .din14(r14tomtree0),
    .din15(r15tomtree0),
    .din16(r16tomtree0),
    .din17(r17tomtree0),
    .din18(r18tomtree0),
    .din19(r19tomtree0),
    .din20(r20tomtree0),
    .din21(r21tomtree0),
    .din22(r22tomtree0),
    .din23(r23tomtree0),
    .din24(r24tomtree0),
    .din25(r25tomtree0),
    .din26(r26tomtree0),
    .din27(r27tomtree0),
    .din28(r28tomtree0),
    .din29(r29tomtree0),
    .din30(r30tomtree0),
    .din31(r31tomtree0),
    .din32(r32tomtree0),
    .din33(r33tomtree0),
    .din34(r34tomtree0),
    .din35(r35tomtree0),
    .din36(r36tomtree0),
    .din37(r37tomtree0),
    .din38(r38tomtree0),
    .din39(r39tomtree0),
    .din40(r40tomtree0),
    .din41(r41tomtree0),
    .din42(r42tomtree0),
    .din43(r43tomtree0),
    .din44(r44tomtree0),
    .din45(r45tomtree0),
    .din46(r46tomtree0),
    .din47(r47tomtree0),
    .din48(r48tomtree0),
    .din49(r49tomtree0),
    .din50(r50tomtree0),
    .din51(r51tomtree0),
    .din52(r52tomtree0),
    .din53(r53tomtree0),
    .din54(r54tomtree0),
    .din55(r55tomtree0),
    .din56(r56tomtree0),
    .din57(r57tomtree0),
    .din58(r58tomtree0),
    .din59(r59tomtree0),
    .din60(r60tomtree0),
    .din61(r61tomtree0),
    .din62(r62tomtree0),
    .din63(r63tomtree0),
    .din64(r64tomtree0),
    .din65(r65tomtree0),
    .din66(r66tomtree0),
    .din67(r67tomtree0),
    .din68(r68tomtree0),
    .din69(r69tomtree0),
    .din70(r70tomtree0),
    .din71(r71tomtree0),
    .din72(r72tomtree0),
    .din73(r73tomtree0),
    .din74(r74tomtree0),
    .din75(r75tomtree0),
    .din76(r76tomtree0),
    .din77(r77tomtree0),
    .din78(r78tomtree0),
    .din79(r79tomtree0),
    .din80(r80tomtree0),
    .din81(r81tomtree0),
    .din82(r82tomtree0),
    .din83(r83tomtree0),
    .din84(r84tomtree0),
    .din85(r85tomtree0),
    .din86(r86tomtree0),
    .din87(r87tomtree0),
    .din88(r88tomtree0),
    .din89(r89tomtree0),
    .din90(r90tomtree0),
    .din91(r91tomtree0),
    .din92(r92tomtree0),
    .din93(r93tomtree0),
    .din94(r94tomtree0),
    .din95(r95tomtree0),
    .din96(r96tomtree0),
    .din97(r97tomtree0),
    .din98(r98tomtree0),
    .din99(r99tomtree0),
    .din100(r100tomtree0),
    .din101(r101tomtree0),
    .din102(r102tomtree0),
    .din103(r103tomtree0),
    .din104(r104tomtree0),
    .din105(r105tomtree0),
    .din106(r106tomtree0),
    .din107(r107tomtree0),
    .din108(r108tomtree0),
    .din109(r109tomtree0),
    .din110(r110tomtree0),
    .din111(r111tomtree0),
    .din112(r112tomtree0),
    .din113(r113tomtree0),
    .din114(r114tomtree0),
    .din115(r115tomtree0),
    .din116(r116tomtree0),
    .din117(r117tomtree0),
    .din118(r118tomtree0),
    .din119(r119tomtree0),
    .din120(r120tomtree0),
    .din121(r121tomtree0),
    .din122(r122tomtree0),
    .din123(r123tomtree0),
    .din124(r124tomtree0),
    .din125(r125tomtree0),
    .din126(r126tomtree0),
    .din127(r127tomtree0),
    .din128(r128tomtree1),
    .din129(r129tomtree1),
    .din130(r130tomtree1),
    .din131(r131tomtree1),
    .din132(r132tomtree1),
    .din133(r133tomtree1),
    .din134(r134tomtree1),
    .din135(r135tomtree1),
    .din136(r136tomtree1),
    .din137(r137tomtree1),
    .din138(r138tomtree1),
    .din139(r139tomtree1),
    .din140(r140tomtree1),
    .din141(r141tomtree1),
    .din142(r142tomtree1),
    .din143(r143tomtree1),
    .din144(r144tomtree1),
    .din145(r145tomtree1),
    .din146(r146tomtree1),
    .din147(r147tomtree1),
    .din148(r148tomtree1),
    .din149(r149tomtree1),
    .din150(r150tomtree1),
    .din151(r151tomtree1),
    .din152(r152tomtree1),
    .din153(r153tomtree1),
    .din154(r154tomtree1),
    .din155(r155tomtree1),
    .din156(r156tomtree1),
    .din157(r157tomtree1),
    .din158(r158tomtree1),
    .din159(r159tomtree1),
    .din160(r160tomtree1),
    .din161(r161tomtree1),
    .din162(r162tomtree1),
    .din163(r163tomtree1),
    .din164(r164tomtree1),
    .din165(r165tomtree1),
    .din166(r166tomtree1),
    .din167(r167tomtree1),
    .din168(r168tomtree1),
    .din169(r169tomtree1),
    .din170(r170tomtree1),
    .din171(r171tomtree1),
    .din172(r172tomtree1),
    .din173(r173tomtree1),
    .din174(r174tomtree1),
    .din175(r175tomtree1),
    .din176(r176tomtree1),
    .din177(r177tomtree1),
    .din178(r178tomtree1),
    .din179(r179tomtree1),
    .din180(r180tomtree1),
    .din181(r181tomtree1),
    .din182(r182tomtree1),
    .din183(r183tomtree1),
    .din184(r184tomtree1),
    .din185(r185tomtree1),
    .din186(r186tomtree1),
    .din187(r187tomtree1),
    .din188(r188tomtree1),
    .din189(r189tomtree1),
    .din190(r190tomtree1),
    .din191(r191tomtree1),
    .din192(r192tomtree1),
    .din193(r193tomtree1),
    .din194(r194tomtree1),
    .din195(r195tomtree1),
    .din196(r196tomtree1),
    .din197(r197tomtree1),
    .din198(r198tomtree1),
    .din199(r199tomtree1),
    .din200(r200tomtree1),
    .din201(r201tomtree1),
    .din202(r202tomtree1),
    .din203(r203tomtree1),
    .din204(r204tomtree1),
    .din205(r205tomtree1),
    .din206(r206tomtree1),
    .din207(r207tomtree1),
    .din208(r208tomtree1),
    .din209(r209tomtree1),
    .din210(r210tomtree1),
    .din211(r211tomtree1),
    .din212(r212tomtree1),
    .din213(r213tomtree1),
    .din214(r214tomtree1),
    .din215(r215tomtree1),
    .din216(r216tomtree1),
    .din217(r217tomtree1),
    .din218(r218tomtree1),
    .din219(r219tomtree1),
    .din220(r220tomtree1),
    .din221(r221tomtree1),
    .din222(r222tomtree1),
    .din223(r223tomtree1),
    .din224(r224tomtree1),
    .din225(r225tomtree1),
    .din226(r226tomtree1),
    .din227(r227tomtree1),
    .din228(r228tomtree1),
    .din229(r229tomtree1),
    .din230(r230tomtree1),
    .din231(r231tomtree1),
    .din232(r232tomtree1),
    .din233(r233tomtree1),
    .din234(r234tomtree1),
    .din235(r235tomtree1),
    .din236(r236tomtree1),
    .din237(r237tomtree1),
    .din238(r238tomtree1),
    .din239(r239tomtree1),
    .din240(r240tomtree1),
    .din241(r241tomtree1),
    .din242(r242tomtree1),
    .din243(r243tomtree1),
    .din244(r244tomtree1),
    .din245(r245tomtree1),
    .din246(r246tomtree1),
    .din247(r247tomtree1),
    .din248(r248tomtree1),
    .din249(r249tomtree1),
    .din250(r250tomtree1),
    .din251(r251tomtree1),
    .din252(r252tomtree1),
    .din253(r253tomtree1),
    .din254(r254tomtree1),
    .din255(r255tomtree1),
    .din256(r256tomtree2),
    .din257(r257tomtree2),
    .din258(r258tomtree2),
    .din259(r259tomtree2),
    .din260(r260tomtree2),
    .din261(r261tomtree2),
    .din262(r262tomtree2),
    .din263(r263tomtree2),
    .din264(r264tomtree2),
    .din265(r265tomtree2),
    .din266(r266tomtree2),
    .din267(r267tomtree2),
    .din268(r268tomtree2),
    .din269(r269tomtree2),
    .din270(r270tomtree2),
    .din271(r271tomtree2),
    .din272(r272tomtree2),
    .din273(r273tomtree2),
    .din274(r274tomtree2),
    .din275(r275tomtree2),
    .din276(r276tomtree2),
    .din277(r277tomtree2),
    .din278(r278tomtree2),
    .din279(r279tomtree2),
    .din280(r280tomtree2),
    .din281(r281tomtree2),
    .din282(r282tomtree2),
    .din283(r283tomtree2),
    .din284(r284tomtree2),
    .din285(r285tomtree2),
    .din286(r286tomtree2),
    .din287(r287tomtree2),
    .din288(r288tomtree2),
    .din289(r289tomtree2),
    .din290(r290tomtree2),
    .din291(r291tomtree2),
    .din292(r292tomtree2),
    .din293(r293tomtree2),
    .din294(r294tomtree2),
    .din295(r295tomtree2),
    .din296(r296tomtree2),
    .din297(r297tomtree2),
    .din298(r298tomtree2),
    .din299(r299tomtree2),
    .din300(r300tomtree2),
    .din301(r301tomtree2),
    .din302(r302tomtree2),
    .din303(r303tomtree2),
    .din304(r304tomtree2),
    .din305(r305tomtree2),
    .din306(r306tomtree2),
    .din307(r307tomtree2),
    .din308(r308tomtree2),
    .din309(r309tomtree2),
    .din310(r310tomtree2),
    .din311(r311tomtree2),
    .din312(r312tomtree2),
    .din313(r313tomtree2),
    .din314(r314tomtree2),
    .din315(r315tomtree2),
    .din316(r316tomtree2),
    .din317(r317tomtree2),
    .din318(r318tomtree2),
    .din319(r319tomtree2),
    .din320(r320tomtree2),
    .din321(r321tomtree2),
    .din322(r322tomtree2),
    .din323(r323tomtree2),
    .din324(r324tomtree2),
    .din325(r325tomtree2),
    .din326(r326tomtree2),
    .din327(r327tomtree2),
    .din328(r328tomtree2),
    .din329(r329tomtree2),
    .din330(r330tomtree2),
    .din331(r331tomtree2),
    .din332(r332tomtree2),
    .din333(r333tomtree2),
    .din334(r334tomtree2),
    .din335(r335tomtree2),
    .din336(r336tomtree2),
    .din337(r337tomtree2),
    .din338(r338tomtree2),
    .din339(r339tomtree2),
    .din340(r340tomtree2),
    .din341(r341tomtree2),
    .din342(r342tomtree2),
    .din343(r343tomtree2),
    .din344(r344tomtree2),
    .din345(r345tomtree2),
    .din346(r346tomtree2),
    .din347(r347tomtree2),
    .din348(r348tomtree2),
    .din349(r349tomtree2),
    .din350(r350tomtree2),
    .din351(r351tomtree2),
    .din352(r352tomtree2),
    .din353(r353tomtree2),
    .din354(r354tomtree2),
    .din355(r355tomtree2),
    .din356(r356tomtree2),
    .din357(r357tomtree2),
    .din358(r358tomtree2),
    .din359(r359tomtree2),
    .din360(r360tomtree2),
    .din361(r361tomtree2),
    .din362(r362tomtree2),
    .din363(r363tomtree2),
    .din364(r364tomtree2),
    .din365(r365tomtree2),
    .din366(r366tomtree2),
    .din367(r367tomtree2),
    .din368(r368tomtree2),
    .din369(r369tomtree2),
    .din370(r370tomtree2),
    .din371(r371tomtree2),
    .din372(r372tomtree2),
    .din373(r373tomtree2),
    .din374(r374tomtree2),
    .din375(r375tomtree2),
    .din376(r376tomtree2),
    .din377(r377tomtree2),
    .din378(r378tomtree2),
    .din379(r379tomtree2),
    .din380(r380tomtree2),
    .din381(r381tomtree2),
    .din382(r382tomtree2),
    .din383(r383tomtree2),
    .din384(r384tomtree3),
    .din385(r385tomtree3),
    .din386(r386tomtree3),
    .din387(r387tomtree3),
    .din388(r388tomtree3),
    .din389(r389tomtree3),
    .din390(r390tomtree3),
    .din391(r391tomtree3),
    .din392(r392tomtree3),
    .din393(r393tomtree3),
    .din394(r394tomtree3),
    .din395(r395tomtree3),
    .din396(r396tomtree3),
    .din397(r397tomtree3),
    .din398(r398tomtree3),
    .din399(r399tomtree3),
    .din400(r400tomtree3),
    .din401(r401tomtree3),
    .din402(r402tomtree3),
    .din403(r403tomtree3),
    .din404(r404tomtree3),
    .din405(r405tomtree3),
    .din406(r406tomtree3),
    .din407(r407tomtree3),
    .din408(r408tomtree3),
    .din409(r409tomtree3),
    .din410(r410tomtree3),
    .din411(r411tomtree3),
    .din412(r412tomtree3),
    .din413(r413tomtree3),
    .din414(r414tomtree3),
    .din415(r415tomtree3),
    .din416(r416tomtree3),
    .din417(r417tomtree3),
    .din418(r418tomtree3),
    .din419(r419tomtree3),
    .din420(r420tomtree3),
    .din421(r421tomtree3),
    .din422(r422tomtree3),
    .din423(r423tomtree3),
    .din424(r424tomtree3),
    .din425(r425tomtree3),
    .din426(r426tomtree3),
    .din427(r427tomtree3),
    .din428(r428tomtree3),
    .din429(r429tomtree3),
    .din430(r430tomtree3),
    .din431(r431tomtree3),
    .din432(r432tomtree3),
    .din433(r433tomtree3),
    .din434(r434tomtree3),
    .din435(r435tomtree3),
    .din436(r436tomtree3),
    .din437(r437tomtree3),
    .din438(r438tomtree3),
    .din439(r439tomtree3),
    .din440(r440tomtree3),
    .din441(r441tomtree3),
    .din442(r442tomtree3),
    .din443(r443tomtree3),
    .din444(r444tomtree3),
    .din445(r445tomtree3),
    .din446(r446tomtree3),
    .din447(r447tomtree3),
    .din448(r448tomtree3),
    .din449(r449tomtree3),
    .din450(r450tomtree3),
    .din451(r451tomtree3),
    .din452(r452tomtree3),
    .din453(r453tomtree3),
    .din454(r454tomtree3),
    .din455(r455tomtree3),
    .din456(r456tomtree3),
    .din457(r457tomtree3),
    .din458(r458tomtree3),
    .din459(r459tomtree3),
    .din460(r460tomtree3),
    .din461(r461tomtree3),
    .din462(r462tomtree3),
    .din463(r463tomtree3),
    .din464(r464tomtree3),
    .din465(r465tomtree3),
    .din466(r466tomtree3),
    .din467(r467tomtree3),
    .din468(r468tomtree3),
    .din469(r469tomtree3),
    .din470(r470tomtree3),
    .din471(r471tomtree3),
    .din472(r472tomtree3),
    .din473(r473tomtree3),
    .din474(r474tomtree3),
    .din475(r475tomtree3),
    .din476(r476tomtree3),
    .din477(r477tomtree3),
    .din478(r478tomtree3),
    .din479(r479tomtree3),
    .din480(r480tomtree3),
    .din481(r481tomtree3),
    .din482(r482tomtree3),
    .din483(r483tomtree3),
    .din484(r484tomtree3),
    .din485(r485tomtree3),
    .din486(r486tomtree3),
    .din487(r487tomtree3),
    .din488(r488tomtree3),
    .din489(r489tomtree3),
    .din490(r490tomtree3),
    .din491(r491tomtree3),
    .din492(r492tomtree3),
    .din493(r493tomtree3),
    .din494(r494tomtree3),
    .din495(r495tomtree3),
    .din496(r496tomtree3),
    .din497(r497tomtree3),
    .din498(r498tomtree3),
    .din499(r499tomtree3),
    .din500(r500tomtree3),
    .din501(r501tomtree3),
    .din502(r502tomtree3),
    .din503(r503tomtree3),
    .din504(r504tomtree3),
    .din505(r505tomtree3),
    .din506(r506tomtree3),
    .din507(r507tomtree3),
    .din508(r508tomtree3),
    .din509(r509tomtree3),
    .din510(r510tomtree3),
    .din511(r511tomtree3),
    .din511(r511tomtree3),
    .din512(r512tomtree4),
    .din513(r513tomtree4),
    .din514(r514tomtree4),
    .din515(r515tomtree4),
    .din516(r516tomtree4),
    .din517(r517tomtree4),
    .din518(r518tomtree4),
    .din519(r519tomtree4),
    .din520(r520tomtree4),
    .din521(r521tomtree4),
    .din522(r522tomtree4),
    .din523(r523tomtree4),
    .din524(r524tomtree4),
    .din525(r525tomtree4),
    .din526(r526tomtree4),
    .din527(r527tomtree4),
    .din528(r528tomtree4),
    .din529(r529tomtree4),
    .din530(r530tomtree4),
    .din531(r531tomtree4),
    .din532(r532tomtree4),
    .din533(r533tomtree4),
    .din534(r534tomtree4),
    .din535(r535tomtree4),
    .din536(r536tomtree4),
    .din537(r537tomtree4),
    .din538(r538tomtree4),
    .din539(r539tomtree4),
    .din540(r540tomtree4),
    .din541(r541tomtree4),
    .din542(r542tomtree4),
    .din543(r543tomtree4),
    .din544(r544tomtree4),
    .din545(r545tomtree4),
    .din546(r546tomtree4),
    .din547(r547tomtree4),
    .din548(r548tomtree4),
    .din549(r549tomtree4),
    .din550(r550tomtree4),
    .din551(r551tomtree4),
    .din552(r552tomtree4),
    .din553(r553tomtree4),
    .din554(r554tomtree4),
    .din555(r555tomtree4),
    .din556(r556tomtree4),
    .din557(r557tomtree4),
    .din558(r558tomtree4),
    .din559(r559tomtree4),
    .din560(r560tomtree4),
    .din561(r561tomtree4),
    .din562(r562tomtree4),
    .din563(r563tomtree4),
    .din564(r564tomtree4),
    .din565(r565tomtree4),
    .din566(r566tomtree4),
    .din567(r567tomtree4),
    .din568(r568tomtree4),
    .din569(r569tomtree4),
    .din570(r570tomtree4),
    .din571(r571tomtree4),
    .din572(r572tomtree4),
    .din573(r573tomtree4),
    .din574(r574tomtree4),
    .din575(r575tomtree4),
    .din576(r576tomtree4),
    .din577(r577tomtree4),
    .din578(r578tomtree4),
    .din579(r579tomtree4),
    .din580(r580tomtree4),
    .din581(r581tomtree4),
    .din582(r582tomtree4),
    .din583(r583tomtree4),
    .din584(r584tomtree4),
    .din585(r585tomtree4),
    .din586(r586tomtree4),
    .din587(r587tomtree4),
    .din588(r588tomtree4),
    .din589(r589tomtree4),
    .din590(r590tomtree4),
    .din591(r591tomtree4),
    .din592(r592tomtree4),
    .din593(r593tomtree4),
    .din594(r594tomtree4),
    .din595(r595tomtree4),
    .din596(r596tomtree4),
    .din597(r597tomtree4),
    .din598(r598tomtree4),
    .din599(r599tomtree4),
    .din600(r600tomtree4),
    .din601(r601tomtree4),
    .din602(r602tomtree4),
    .din603(r603tomtree4),
    .din604(r604tomtree4),
    .din605(r605tomtree4),
    .din606(r606tomtree4),
    .din607(r607tomtree4),
    .din608(r608tomtree4),
    .din609(r609tomtree4),
    .din610(r610tomtree4),
    .din611(r611tomtree4),
    .din612(r612tomtree4),
    .din613(r613tomtree4),
    .din614(r614tomtree4),
    .din615(r615tomtree4),
    .din616(r616tomtree4),
    .din617(r617tomtree4),
    .din618(r618tomtree4),
    .din619(r619tomtree4),
    .din620(r620tomtree4),
    .din621(r621tomtree4),
    .din622(r622tomtree4),
    .din623(r623tomtree4),
    .din624(r624tomtree4),
    .din625(r625tomtree4),
    .din626(r626tomtree4),
    .din627(r627tomtree4),
    .din628(r628tomtree4),
    .din629(r629tomtree4),
    .din630(r630tomtree4),
    .din631(r631tomtree4),
    .din632(r632tomtree4),
    .din633(r633tomtree4),
    .din634(r634tomtree4),
    .din635(r635tomtree4),
    .din636(r636tomtree4),
    .din637(r637tomtree4),
    .din638(r638tomtree4),
    .din639(r639tomtree4),
    .din640(r640tomtree5),
    .din641(r641tomtree5),
    .din642(r642tomtree5),
    .din643(r643tomtree5),
    .din644(r644tomtree5),
    .din645(r645tomtree5),
    .din646(r646tomtree5),
    .din647(r647tomtree5),
    .din648(r648tomtree5),
    .din649(r649tomtree5),
    .din650(r650tomtree5),
    .din651(r651tomtree5),
    .din652(r652tomtree5),
    .din653(r653tomtree5),
    .din654(r654tomtree5),
    .din655(r655tomtree5),
    .din656(r656tomtree5),
    .din657(r657tomtree5),
    .din658(r658tomtree5),
    .din659(r659tomtree5),
    .din660(r660tomtree5),
    .din661(r661tomtree5),
    .din662(r662tomtree5),
    .din663(r663tomtree5),
    .din664(r664tomtree5),
    .din665(r665tomtree5),
    .din666(r666tomtree5),
    .din667(r667tomtree5),
    .din668(r668tomtree5),
    .din669(r669tomtree5),
    .din670(r670tomtree5),
    .din671(r671tomtree5),
    .din672(r672tomtree5),
    .din673(r673tomtree5),
    .din674(r674tomtree5),
    .din675(r675tomtree5),
    .din676(r676tomtree5),
    .din677(r677tomtree5),
    .din678(r678tomtree5),
    .din679(r679tomtree5),
    .din680(r680tomtree5),
    .din681(r681tomtree5),
    .din682(r682tomtree5),
    .din683(r683tomtree5),
    .din684(r684tomtree5),
    .din685(r685tomtree5),
    .din686(r686tomtree5),
    .din687(r687tomtree5),
    .din688(r688tomtree5),
    .din689(r689tomtree5),
    .din690(r690tomtree5),
    .din691(r691tomtree5),
    .din692(r692tomtree5),
    .din693(r693tomtree5),
    .din694(r694tomtree5),
    .din695(r695tomtree5),
    .din696(r696tomtree5),
    .din697(r697tomtree5),
    .din698(r698tomtree5),
    .din699(r699tomtree5),
    .din700(r700tomtree5),
    .din701(r701tomtree5),
    .din702(r702tomtree5),
    .din703(r703tomtree5),
    .din704(r704tomtree5),
    .din705(r705tomtree5),
    .din706(r706tomtree5),
    .din707(r707tomtree5),
    .din708(r708tomtree5),
    .din709(r709tomtree5),
    .din710(r710tomtree5),
    .din711(r711tomtree5),
    .din712(r712tomtree5),
    .din713(r713tomtree5),
    .din714(r714tomtree5),
    .din715(r715tomtree5),
    .din716(r716tomtree5),
    .din717(r717tomtree5),
    .din718(r718tomtree5),
    .din719(r719tomtree5),
    .din720(r720tomtree5),
    .din721(r721tomtree5),
    .din722(r722tomtree5),
    .din723(r723tomtree5),
    .din724(r724tomtree5),
    .din725(r725tomtree5),
    .din726(r726tomtree5),
    .din727(r727tomtree5),
    .din728(r728tomtree5),
    .din729(r729tomtree5),
    .din730(r730tomtree5),
    .din731(r731tomtree5),
    .din732(r732tomtree5),
    .din733(r733tomtree5),
    .din734(r734tomtree5),
    .din735(r735tomtree5),
    .din736(r736tomtree5),
    .din737(r737tomtree5),
    .din738(r738tomtree5),
    .din739(r739tomtree5),
    .din740(r740tomtree5),
    .din741(r741tomtree5),
    .din742(r742tomtree5),
    .din743(r743tomtree5),
    .din744(r744tomtree5),
    .din745(r745tomtree5),
    .din746(r746tomtree5),
    .din747(r747tomtree5),
    .din748(r748tomtree5),
    .din749(r749tomtree5),
    .din750(r750tomtree5),
    .din751(r751tomtree5),
    .din752(r752tomtree5),
    .din753(r753tomtree5),
    .din754(r754tomtree5),
    .din755(r755tomtree5),
    .din756(r756tomtree5),
    .din757(r757tomtree5),
    .din758(r758tomtree5),
    .din759(r759tomtree5),
    .din760(r760tomtree5),
    .din761(r761tomtree5),
    .din762(r762tomtree5),
    .din763(r763tomtree5),
    .din764(r764tomtree5),
    .din765(r765tomtree5),
    .din766(r766tomtree5),
    .din767(r767tomtree5),
    .din768(r768tomtree6),
    .din769(r769tomtree6),
    .din770(r770tomtree6),
    .din771(r771tomtree6),
    .din772(r772tomtree6),
    .din773(r773tomtree6),
    .din774(r774tomtree6),
    .din775(r775tomtree6),
    .din776(r776tomtree6),
    .din777(r777tomtree6),
    .din778(r778tomtree6),
    .din779(r779tomtree6),
    .din780(r780tomtree6),
    .din781(r781tomtree6),
    .din782(r782tomtree6),
    .din783(r783tomtree6),
    .din784(r784tomtree6),
    .din785(r785tomtree6),
    .din786(r786tomtree6),
    .din787(r787tomtree6),
    .din788(r788tomtree6),
    .din789(r789tomtree6),
    .din790(r790tomtree6),
    .din791(r791tomtree6),
    .din792(r792tomtree6),
    .din793(r793tomtree6),
    .din794(r794tomtree6),
    .din795(r795tomtree6),
    .din796(r796tomtree6),
    .din797(r797tomtree6),
    .din798(r798tomtree6),
    .din799(r799tomtree6),
    .din800(r800tomtree6),
    .din801(r801tomtree6),
    .din802(r802tomtree6),
    .din803(r803tomtree6),
    .din804(r804tomtree6),
    .din805(r805tomtree6),
    .din806(r806tomtree6),
    .din807(r807tomtree6),
    .din808(r808tomtree6),
    .din809(r809tomtree6),
    .din810(r810tomtree6),
    .din811(r811tomtree6),
    .din812(r812tomtree6),
    .din813(r813tomtree6),
    .din814(r814tomtree6),
    .din815(r815tomtree6),
    .din816(r816tomtree6),
    .din817(r817tomtree6),
    .din818(r818tomtree6),
    .din819(r819tomtree6),
    .din820(r820tomtree6),
    .din821(r821tomtree6),
    .din822(r822tomtree6),
    .din823(r823tomtree6),
    .din824(r824tomtree6),
    .din825(r825tomtree6),
    .din826(r826tomtree6),
    .din827(r827tomtree6),
    .din828(r828tomtree6),
    .din829(r829tomtree6),
    .din830(r830tomtree6),
    .din831(r831tomtree6),
    .din832(r832tomtree6),
    .din833(r833tomtree6),
    .din834(r834tomtree6),
    .din835(r835tomtree6),
    .din836(r836tomtree6),
    .din837(r837tomtree6),
    .din838(r838tomtree6),
    .din839(r839tomtree6),
    .din840(r840tomtree6),
    .din841(r841tomtree6),
    .din842(r842tomtree6),
    .din843(r843tomtree6),
    .din844(r844tomtree6),
    .din845(r845tomtree6),
    .din846(r846tomtree6),
    .din847(r847tomtree6),
    .din848(r848tomtree6),
    .din849(r849tomtree6),
    .din850(r850tomtree6),
    .din851(r851tomtree6),
    .din852(r852tomtree6),
    .din853(r853tomtree6),
    .din854(r854tomtree6),
    .din855(r855tomtree6),
    .din856(r856tomtree6),
    .din857(r857tomtree6),
    .din858(r858tomtree6),
    .din859(r859tomtree6),
    .din860(r860tomtree6),
    .din861(r861tomtree6),
    .din862(r862tomtree6),
    .din863(r863tomtree6),
    .din864(r864tomtree6),
    .din865(r865tomtree6),
    .din866(r866tomtree6),
    .din867(r867tomtree6),
    .din868(r868tomtree6),
    .din869(r869tomtree6),
    .din870(r870tomtree6),
    .din871(r871tomtree6),
    .din872(r872tomtree6),
    .din873(r873tomtree6),
    .din874(r874tomtree6),
    .din875(r875tomtree6),
    .din876(r876tomtree6),
    .din877(r877tomtree6),
    .din878(r878tomtree6),
    .din879(r879tomtree6),
    .din880(r880tomtree6),
    .din881(r881tomtree6),
    .din882(r882tomtree6),
    .din883(r883tomtree6),
    .din884(r884tomtree6),
    .din885(r885tomtree6),
    .din886(r886tomtree6),
    .din887(r887tomtree6),
    .din888(r888tomtree6),
    .din889(r889tomtree6),
    .din890(r890tomtree6),
    .din891(r891tomtree6),
    .din892(r892tomtree6),
    .din893(r893tomtree6),
    .din894(r894tomtree6),
    .din895(r895tomtree6),
    .din896(r896tomtree7),
    .din897(r897tomtree7),
    .din898(r898tomtree7),
    .din899(r899tomtree7),
    .din900(r900tomtree7),
    .din901(r901tomtree7),
    .din902(r902tomtree7),
    .din903(r903tomtree7),
    .din904(r904tomtree7),
    .din905(r905tomtree7),
    .din906(r906tomtree7),
    .din907(r907tomtree7),
    .din908(r908tomtree7),
    .din909(r909tomtree7),
    .din910(r910tomtree7),
    .din911(r911tomtree7),
    .din912(r912tomtree7),
    .din913(r913tomtree7),
    .din914(r914tomtree7),
    .din915(r915tomtree7),
    .din916(r916tomtree7),
    .din917(r917tomtree7),
    .din918(r918tomtree7),
    .din919(r919tomtree7),
    .din920(r920tomtree7),
    .din921(r921tomtree7),
    .din922(r922tomtree7),
    .din923(r923tomtree7),
    .din924(r924tomtree7),
    .din925(r925tomtree7),
    .din926(r926tomtree7),
    .din927(r927tomtree7),
    .din928(r928tomtree7),
    .din929(r929tomtree7),
    .din930(r930tomtree7),
    .din931(r931tomtree7),
    .din932(r932tomtree7),
    .din933(r933tomtree7),
    .din934(r934tomtree7),
    .din935(r935tomtree7),
    .din936(r936tomtree7),
    .din937(r937tomtree7),
    .din938(r938tomtree7),
    .din939(r939tomtree7),
    .din940(r940tomtree7),
    .din941(r941tomtree7),
    .din942(r942tomtree7),
    .din943(r943tomtree7),
    .din944(r944tomtree7),
    .din945(r945tomtree7),
    .din946(r946tomtree7),
    .din947(r947tomtree7),
    .din948(r948tomtree7),
    .din949(r949tomtree7),
    .din950(r950tomtree7),
    .din951(r951tomtree7),
    .din952(r952tomtree7),
    .din953(r953tomtree7),
    .din954(r954tomtree7),
    .din955(r955tomtree7),
    .din956(r956tomtree7),
    .din957(r957tomtree7),
    .din958(r958tomtree7),
    .din959(r959tomtree7),
    .din960(r960tomtree7),
    .din961(r961tomtree7),
    .din962(r962tomtree7),
    .din963(r963tomtree7),
    .din964(r964tomtree7),
    .din965(r965tomtree7),
    .din966(r966tomtree7),
    .din967(r967tomtree7),
    .din968(r968tomtree7),
    .din969(r969tomtree7),
    .din970(r970tomtree7),
    .din971(r971tomtree7),
    .din972(r972tomtree7),
    .din973(r973tomtree7),
    .din974(r974tomtree7),
    .din975(r975tomtree7),
    .din976(r976tomtree7),
    .din977(r977tomtree7),
    .din978(r978tomtree7),
    .din979(r979tomtree7),
    .din980(r980tomtree7),
    .din981(r981tomtree7),
    .din982(r982tomtree7),
    .din983(r983tomtree7),
    .din984(r984tomtree7),
    .din985(r985tomtree7),
    .din986(r986tomtree7),
    .din987(r987tomtree7),
    .din988(r988tomtree7),
    .din989(r989tomtree7),
    .din990(r990tomtree7),
    .din991(r991tomtree7),
    .din992(r992tomtree7),
    .din993(r993tomtree7),
    .din994(r994tomtree7),
    .din995(r995tomtree7),
    .din996(r996tomtree7),
    .din997(r997tomtree7),
    .din998(r998tomtree7),
    .din999(r999tomtree7),
    .din1000(r1000tomtree7),
    .din1001(r1001tomtree7),
    .din1002(r1002tomtree7),
    .din1003(r1003tomtree7),
    .din1004(r1004tomtree7),
    .din1005(r1005tomtree7),
    .din1006(r1006tomtree7),
    .din1007(r1007tomtree7),
    .din1008(r1008tomtree7),
    .din1009(r1009tomtree7),
    .din1010(r1010tomtree7),
    .din1011(r1011tomtree7),
    .din1012(r1012tomtree7),
    .din1013(r1013tomtree7),
    .din1014(r1014tomtree7),
    .din1015(r1015tomtree7),
    .din1016(r1016tomtree7),
    .din1017(r1017tomtree7),
    .din1018(r1018tomtree7),
    .din1019(r1019tomtree7),
    .din1020(r1020tomtree7),
    .din1021(r1021tomtree7),
    .din1022(r1022tomtree7),
    .din1023(r1023tomtree7),
    .sel(cntout),
    .indx(indx)
  );

  counter_out #(.INCR(1), .CNT_WIDTH($clog2(BATCH_SIZE))) CntOut(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntouten),
    .cnt(cntout)
  );

  counter_addr #(.INCR(ADDR_INCR_PORTB), .ADDR_WIDTH(ADDR_WIDTH_PORTB)) CntAddrB(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntaddrben),
    .cnt(addrbw)
  );
  
  //bram output port
  assign clkb = clk;
  assign rstb = ~rst_n;
  assign enb = enbw;
  assign addrb = addrbw;
  assign dinb = indx;
  assign web = webw;
  
endmodule