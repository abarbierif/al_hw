`timescale 1ns / 1ps

module margin_sampling10(
  input  wire clk,
  input  wire rst_n,
  // *** CONTROL AND STATUS PORT ***
  output wire ready,
  input  wire start,
  // *** DATA INPUT PORT ***
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA CLK" *)  output wire clka,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA RST" *)  output wire rsta,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA EN" *)   output wire ena,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA ADDR" *) output wire [31:0] addra,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA DIN" *)  output wire [255:0] dina,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA WE" *)   output wire [31:0] wea,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTA DOUT" *) input  wire [255:0] douta,
  // *** DATA OUTPUT PORT ***
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB CLK" *)  output wire clkb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB RST" *)  output wire rstb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB EN" *)   output wire enb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB ADDR" *) output wire [31:0] addrb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB DIN" *)  output wire [31:0] dinb,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB WE" *)   output wire [3:0] web,
  (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 BRAM_PORTB DOUT" *) input  wire [31:0] doutb
);
  
  //local parameters
  localparam DATA_WIDTH = 16;
  localparam BATCH_SIZE = 512;
  localparam MAX_DATA_LENGTH = 10*BATCH_SIZE;
  localparam DATA_LENGTH = 5120;
  localparam ADDR_WIDTH_PORTA = 32;
  localparam ADDR_INCR_PORTA = 32;
  localparam ADDR_WIDTH_PORTB = 32;
  localparam ADDR_INCR_PORTB = 4;
  localparam N_REGISTERS = 64;
  localparam N_REGISTERSBANKS = 8;
  localparam INDX_WIDTH = $clog2(MAX_DATA_LENGTH);
  localparam ADDR_WIDTH = $clog2(N_REGISTERS);
  localparam MARGIN_PIPELINE_DEPTH = 7;
  
  //wires
  wire startrising;
  
  wire [DATA_WIDTH-1:0] din0, din1, din2, din3, din4, din5, din6, din7, din8, din9;
  wire [DATA_WIDTH-1:0] rdin0, rdin1, rdin2, rdin3, rdin4, rdin5, rdin6, rdin7, rdin8, rdin9;
  wire [DATA_WIDTH-1:0] mrgn;
  
  wire trigmax;
  wire rtrigmax;
  wire enaw;
  wire [31:0] weaw;
  wire enbw;
  wire [3:0] webw;
  wire cntaddraen;
  wire mrgnpipelineen;
  wire cntindxen;  
  wire cntren;
  wire cntrben;
  wire rsrc;  
  wire rbsrc;
  wire decrsrc;
  wire decrbsrc;
  wire mrgnsrc; 
  wire trigmtree;
  wire cntouten;
  wire cntaddrben;
  
  wire [ADDR_WIDTH_PORTA-1:0] addraw;
  wire [ADDR_WIDTH_PORTB-1:0] addrbw;
  wire [INDX_WIDTH-1:0] mrgnindx;
  wire [INDX_WIDTH-1:0] indx;
  wire [$clog2(N_REGISTERS)-1:0] cntr;
  wire [$clog2(N_REGISTERS)-1:0] rcntr;
  wire [$clog2(N_REGISTERSBANKS)-1:0] cntrb; //cntrb0, cntrb1, cntrb2, cntrb3, cntrb4, cntrb5, cntrb6, cntrb7;
  wire [$clog2(N_REGISTERSBANKS)-1:0] rcntrb;
  wire [$clog2(N_REGISTERSBANKS)-1:0] rrcntrb;
  wire [$clog2(N_REGISTERS)-1:0] decrsrcmuxout;
  wire [$clog2(N_REGISTERSBANKS)-1:0] decrbsrcmuxout;
  wire [N_REGISTERS-1:0] decr;
  wire [N_REGISTERSBANKS-1:0] decrb; //decrb0, decrb1, decrb2, decrb3, decrb4, decrb5, decrb6, decrb7;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] mrgnsrcmuxout;
  wire [N_REGISTERS-1:0] rsrcmuxout;
  wire [N_REGISTERSBANKS-1:0] rbsrcmuxout; //rbsrcmuxout0, rbsrcmuxout1, rbsrcmuxout2, rbsrcmuxout3, rbsrcmuxout4, rbsrcmuxout5, rbsrcmuxout6, rbsrcmuxout7;
  
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] r0tomtree0, r1tomtree0, r2tomtree0, r3tomtree0, r4tomtree0, r5tomtree0,
  r6tomtree0, r7tomtree0, r8tomtree0, r9tomtree0, r10tomtree0, r11tomtree0, r12tomtree0, r13tomtree0, r14tomtree0, r15tomtree0,
  r16tomtree0, r17tomtree0, r18tomtree0, r19tomtree0, r20tomtree0, r21tomtree0, r22tomtree0, r23tomtree0, r24tomtree0, r25tomtree0,
  r26tomtree0, r27tomtree0, r28tomtree0, r29tomtree0, r30tomtree0, r31tomtree0, r32tomtree0, r33tomtree0, r34tomtree0, r35tomtree0,
  r36tomtree0, r37tomtree0, r38tomtree0, r39tomtree0, r40tomtree0, r41tomtree0, r42tomtree0, r43tomtree0, r44tomtree0, r45tomtree0,
  r46tomtree0, r47tomtree0, r48tomtree0, r49tomtree0, r50tomtree0, r51tomtree0, r52tomtree0, r53tomtree0, r54tomtree0, r55tomtree0,
  r56tomtree0, r57tomtree0, r58tomtree0, r59tomtree0, r60tomtree0, r61tomtree0, r62tomtree0, r63tomtree0, r64tomtree1, r65tomtree1,
  r66tomtree1, r67tomtree1, r68tomtree1, r69tomtree1, r70tomtree1, r71tomtree1, r72tomtree1, r73tomtree1, r74tomtree1, r75tomtree1,
  r76tomtree1, r77tomtree1, r78tomtree1, r79tomtree1, r80tomtree1, r81tomtree1, r82tomtree1, r83tomtree1, r84tomtree1, r85tomtree1,
  r86tomtree1, r87tomtree1, r88tomtree1, r89tomtree1, r90tomtree1, r91tomtree1, r92tomtree1, r93tomtree1, r94tomtree1, r95tomtree1,
  r96tomtree1, r97tomtree1, r98tomtree1, r99tomtree1, r100tomtree1, r101tomtree1, r102tomtree1, r103tomtree1, r104tomtree1, r105tomtree1,
  r106tomtree1, r107tomtree1, r108tomtree1, r109tomtree1, r110tomtree1, r111tomtree1, r112tomtree1, r113tomtree1, r114tomtree1, r115tomtree1,
  r116tomtree1, r117tomtree1, r118tomtree1, r119tomtree1, r120tomtree1, r121tomtree1, r122tomtree1, r123tomtree1, r124tomtree1, r125tomtree1,
  r126tomtree1, r127tomtree1, r128tomtree2, r129tomtree2, r130tomtree2, r131tomtree2, r132tomtree2, r133tomtree2, r134tomtree2, r135tomtree2,
  r136tomtree2, r137tomtree2, r138tomtree2, r139tomtree2, r140tomtree2, r141tomtree2, r142tomtree2, r143tomtree2, r144tomtree2, r145tomtree2,
  r146tomtree2, r147tomtree2, r148tomtree2, r149tomtree2, r150tomtree2, r151tomtree2, r152tomtree2, r153tomtree2, r154tomtree2, r155tomtree2,
  r156tomtree2, r157tomtree2, r158tomtree2, r159tomtree2, r160tomtree2, r161tomtree2, r162tomtree2, r163tomtree2, r164tomtree2, r165tomtree2,
  r166tomtree2, r167tomtree2, r168tomtree2, r169tomtree2, r170tomtree2, r171tomtree2, r172tomtree2, r173tomtree2, r174tomtree2, r175tomtree2,
  r176tomtree2, r177tomtree2, r178tomtree2, r179tomtree2, r180tomtree2, r181tomtree2, r182tomtree2, r183tomtree2, r184tomtree2, r185tomtree2,
  r186tomtree2, r187tomtree2, r188tomtree2, r189tomtree2, r190tomtree2, r191tomtree2, r192tomtree3, r193tomtree3, r194tomtree3, r195tomtree3,
  r196tomtree3, r197tomtree3, r198tomtree3, r199tomtree3, r200tomtree3, r201tomtree3, r202tomtree3, r203tomtree3, r204tomtree3, r205tomtree3,
  r206tomtree3, r207tomtree3, r208tomtree3, r209tomtree3, r210tomtree3, r211tomtree3, r212tomtree3, r213tomtree3, r214tomtree3, r215tomtree3,
  r216tomtree3, r217tomtree3, r218tomtree3, r219tomtree3, r220tomtree3, r221tomtree3, r222tomtree3, r223tomtree3, r224tomtree3, r225tomtree3,
  r226tomtree3, r227tomtree3, r228tomtree3, r229tomtree3, r230tomtree3, r231tomtree3, r232tomtree3, r233tomtree3, r234tomtree3, r235tomtree3,
  r236tomtree3, r237tomtree3, r238tomtree3, r239tomtree3, r240tomtree3, r241tomtree3, r242tomtree3, r243tomtree3, r244tomtree3, r245tomtree3,
  r246tomtree3, r247tomtree3, r248tomtree3, r249tomtree3, r250tomtree3, r251tomtree3, r252tomtree3, r253tomtree3, r254tomtree3, r255tomtree3,
  r256tomtree4, r257tomtree4, r258tomtree4, r259tomtree4, r260tomtree4, r261tomtree4, r262tomtree4, r263tomtree4, r264tomtree4, r265tomtree4,
  r266tomtree4, r267tomtree4, r268tomtree4, r269tomtree4, r270tomtree4, r271tomtree4, r272tomtree4, r273tomtree4, r274tomtree4, r275tomtree4,
  r276tomtree4, r277tomtree4, r278tomtree4, r279tomtree4, r280tomtree4, r281tomtree4, r282tomtree4, r283tomtree4, r284tomtree4, r285tomtree4,
  r286tomtree4, r287tomtree4, r288tomtree4, r289tomtree4, r290tomtree4, r291tomtree4, r292tomtree4, r293tomtree4, r294tomtree4, r295tomtree4,
  r296tomtree4, r297tomtree4, r298tomtree4, r299tomtree4, r300tomtree4, r301tomtree4, r302tomtree4, r303tomtree4, r304tomtree4, r305tomtree4,
  r306tomtree4, r307tomtree4, r308tomtree4, r309tomtree4, r310tomtree4, r311tomtree4, r312tomtree4, r313tomtree4, r314tomtree4, r315tomtree4,
  r316tomtree4, r317tomtree4, r318tomtree4, r319tomtree4, r320tomtree5, r321tomtree5, r322tomtree5, r323tomtree5, r324tomtree5, r325tomtree5,
  r326tomtree5, r327tomtree5, r328tomtree5, r329tomtree5, r330tomtree5, r331tomtree5, r332tomtree5, r333tomtree5, r334tomtree5, r335tomtree5,
  r336tomtree5, r337tomtree5, r338tomtree5, r339tomtree5, r340tomtree5, r341tomtree5, r342tomtree5, r343tomtree5, r344tomtree5, r345tomtree5,
  r346tomtree5, r347tomtree5, r348tomtree5, r349tomtree5, r350tomtree5, r351tomtree5, r352tomtree5, r353tomtree5, r354tomtree5, r355tomtree5,
  r356tomtree5, r357tomtree5, r358tomtree5, r359tomtree5, r360tomtree5, r361tomtree5, r362tomtree5, r363tomtree5, r364tomtree5, r365tomtree5,
  r366tomtree5, r367tomtree5, r368tomtree5, r369tomtree5, r370tomtree5, r371tomtree5, r372tomtree5, r373tomtree5, r374tomtree5, r375tomtree5,
  r376tomtree5, r377tomtree5, r378tomtree5, r379tomtree5, r380tomtree5, r381tomtree5, r382tomtree5, r383tomtree5, r384tomtree6, r385tomtree6,
  r386tomtree6, r387tomtree6, r388tomtree6, r389tomtree6, r390tomtree6, r391tomtree6, r392tomtree6, r393tomtree6, r394tomtree6, r395tomtree6,
  r396tomtree6, r397tomtree6, r398tomtree6, r399tomtree6, r400tomtree6, r401tomtree6, r402tomtree6, r403tomtree6, r404tomtree6, r405tomtree6,
  r406tomtree6, r407tomtree6, r408tomtree6, r409tomtree6, r410tomtree6, r411tomtree6, r412tomtree6, r413tomtree6, r414tomtree6, r415tomtree6,
  r416tomtree6, r417tomtree6, r418tomtree6, r419tomtree6, r420tomtree6, r421tomtree6, r422tomtree6, r423tomtree6, r424tomtree6, r425tomtree6,
  r426tomtree6, r427tomtree6, r428tomtree6, r429tomtree6, r430tomtree6, r431tomtree6, r432tomtree6, r433tomtree6, r434tomtree6, r435tomtree6,
  r436tomtree6, r437tomtree6, r438tomtree6, r439tomtree6, r440tomtree6, r441tomtree6, r442tomtree6, r443tomtree6, r444tomtree6, r445tomtree6,
  r446tomtree6, r447tomtree6, r448tomtree7, r449tomtree7, r450tomtree7, r451tomtree7, r452tomtree7, r453tomtree7, r454tomtree7, r455tomtree7,
  r456tomtree7, r457tomtree7, r458tomtree7, r459tomtree7, r460tomtree7, r461tomtree7, r462tomtree7, r463tomtree7, r464tomtree7, r465tomtree7,
  r466tomtree7, r467tomtree7, r468tomtree7, r469tomtree7, r470tomtree7, r471tomtree7, r472tomtree7, r473tomtree7, r474tomtree7, r475tomtree7,
  r476tomtree7, r477tomtree7, r478tomtree7, r479tomtree7, r480tomtree7, r481tomtree7, r482tomtree7, r483tomtree7, r484tomtree7, r485tomtree7,
  r486tomtree7, r487tomtree7, r488tomtree7, r489tomtree7, r490tomtree7, r491tomtree7, r492tomtree7, r493tomtree7, r494tomtree7, r495tomtree7,
  r496tomtree7, r497tomtree7, r498tomtree7, r499tomtree7, r500tomtree7, r501tomtree7, r502tomtree7, r503tomtree7, r504tomtree7, r505tomtree7,
  r506tomtree7, r507tomtree7, r508tomtree7, r509tomtree7, r510tomtree7, r511tomtree7;
  
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] mtree0tomaxsrcmux, mtree1tomaxsrcmux, mtree2tomaxsrcmux, 
  mtree3tomaxsrcmux, mtree4tomaxsrcmux, mtree5tomaxsrcmux, mtree6tomaxsrcmux, mtree7tomaxsrcmux;
  
  wire [N_REGISTERSBANKS-1:0] trigmtreesrcmuxout;
  wire [N_REGISTERSBANKS-1:0] trigmtreeold;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] maxsrcmuxtocmp;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] mrgncmp;
  wire [(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)-1:0] rmrgncmp;
  wire [$clog2(N_REGISTERS)-1:0] rcmp;
  wire [$clog2(N_REGISTERS)-1:0] rrcmp; 
  wire [$clog2(BATCH_SIZE)-1:0] cntout;
  
  //start rising
  reg startold;
  always @(posedge clk) begin
    startold <= start;
  end
  assign startrising = !startold && start;
  
  controller #(.DATA_LENGTH(DATA_LENGTH), .MARGIN_PIPELINE_DEPTH(MARGIN_PIPELINE_DEPTH), .N_REGISTERS(N_REGISTERS), .BATCH_SIZE(BATCH_SIZE), .N_REGISTERSBANKS(N_REGISTERSBANKS)) Cntr(
    .clk(clk),
    .rst_n(rst_n),
    .Start(startrising),
    .MTreeSrc(rtrigmax),
    .Ready(ready),
    .EnA(enaw),
    .WeA(weaw),
    .EnB(enbw),
    .WeB(webw),
    .CntAddrAEn(cntaddraen),
    .MrgnPipelineEn(mrgnpipelineen),
    .CntIndxEn(cntindxen),
    .CntREn(cntren),
    .CntRBEn(cntrben),
    .RSrc(rsrc),
    .RBSrc(rbsrc),
    .DecRSrc(decrsrc),
    .DecRBSrc(decrbsrc),
    .MrgnSrc(mrgnsrc),
    .TrigMTree(trigmtree),
    .CntOutEn(cntouten),
    .CntAddrBEn(cntaddrben)
  );

  //bram input port
  assign clka = clk;
  assign rsta = ~rst_n;
  assign ena = enaw;
  assign addra = addraw;
  assign dina = 0;
  assign wea = weaw;
  
  counter_addr #(.INCR(ADDR_INCR_PORTA), .ADDR_WIDTH(ADDR_WIDTH_PORTA)) CntAddrA(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntaddraen),
    .cnt(addraw)
  );
  
  assign din0 = douta[15:0];
  assign din1 = douta[31:16];
  assign din2 = douta[47:32];
  assign din3 = douta[63:48];
  assign din4 = douta[79:64];
  assign din5 = douta[95:80];
  assign din6 = douta[111:96];
  assign din7 = douta[127:112];
  assign din8 = douta[143:128];
  assign din9 = douta[159:144];
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn0(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din0),
    .dout(rdin0)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn1(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din1),
    .dout(rdin1)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn2(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din2),
    .dout(rdin2)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn3(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din3),
    .dout(rdin3)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn4(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din4),
    .dout(rdin4)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn5(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din5),
    .dout(rdin5)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn6(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din6),
    .dout(rdin6)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn7(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din7),
    .dout(rdin7)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn8(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din8),
    .dout(rdin8)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH)) RIn9(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(din9),
    .dout(rdin9)
  );
  
  margin_pipeline10 #(.DATA_WIDTH(DATA_WIDTH)) MrgnPipeline(
    .clk(clk),
    .rst_n(rst_n),
    .en(mrgnpipelineen),
    .din0(rdin0),
    .din1(rdin1),
    .din2(rdin2),
    .din3(rdin3),
    .din4(rdin4),
    .din5(rdin5),
    .din6(rdin6),
    .din7(rdin7),
    .din8(rdin8),
    .din9(rdin9),
    .margin(mrgn)
  );
  
  counter_indx #(.INCR(1), .CNT_WIDTH(INDX_WIDTH)) CntIndx(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntindxen),
    .cnt(mrgnindx)
  );
  
  counter_r #(.MAX_CNT(N_REGISTERS), .INCR(1), .N_REGISTERSBANKS(N_REGISTERSBANKS)) CntR(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntren),
    .cnt(cntr)
  );
  
  register #(.DATA_WIDTH($clog2(N_REGISTERS))) RCntR(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(cntr),
    .dout(rcntr)
  );

  mux2 #(.DATA_WIDTH($clog2(N_REGISTERS))) DecRSrcMux(
    .din0(rcntr), 
    .din1(rrcmp), 
    .sel(decrsrc), 
    .dout(decrsrcmuxout)
  );

  decoder #(.IN_WIDTH($clog2(N_REGISTERS))) DecR(
    .din(decrsrcmuxout), 
    .dout(decr)
  );
  
  counter_rb #(.MAX_CNT(N_REGISTERSBANKS), .INCR(1)) CntRB(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntrben),
    .cnt(cntrb)
  );
  
  register #(.DATA_WIDTH($clog2(N_REGISTERSBANKS))) RCntRB(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(cntrb),
    .dout(rcntrb)
  );
  
  register #(.DATA_WIDTH($clog2(N_REGISTERSBANKS))) RRCntRB(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(rcntrb),
    .dout(rrcntrb)
  );
  
  mux2 #(.DATA_WIDTH($clog2(N_REGISTERSBANKS))) DecRBSrcMux(
    .din0(rcntrb), 
    .din1(rrcntrb), 
    .sel(decrbsrc), 
    .dout(decrbsrcmuxout)
  );

  decoder #(.IN_WIDTH($clog2(N_REGISTERSBANKS))) DecRB(
    .din(decrbsrcmuxout), 
    .dout(decrb)
  );

  mux2 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) MrgnSrcMux(
    .din0(rmrgncmp), 
    .din1({rcntr,mrgnindx,mrgn}), 
    .sel(!mrgnsrc), 
    .dout(mrgnsrcmuxout)
  );

  mux2 #(.DATA_WIDTH(N_REGISTERS)) RSrcMux(
    .din0('b0), 
    .din1(decr), 
    .sel(rsrc), 
    .dout(rsrcmuxout)
  );
  
  mux2 #(.DATA_WIDTH(N_REGISTERSBANKS)) RBSrcMux(
    .din0('b0), 
    .din1(decrb), 
    .sel(rbsrc), 
    .dout(rbsrcmuxout)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_0(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[0]),
    .din(mrgnsrcmuxout),
    .dout0(r0tomtree0),
    .dout1(r1tomtree0),
    .dout2(r2tomtree0),
    .dout3(r3tomtree0),
    .dout4(r4tomtree0),
    .dout5(r5tomtree0),
    .dout6(r6tomtree0),
    .dout7(r7tomtree0),
    .dout8(r8tomtree0),
    .dout9(r9tomtree0),
    .dout10(r10tomtree0),
    .dout11(r11tomtree0),
    .dout12(r12tomtree0),
    .dout13(r13tomtree0),
    .dout14(r14tomtree0),
    .dout15(r15tomtree0),
    .dout16(r16tomtree0),
    .dout17(r17tomtree0),
    .dout18(r18tomtree0),
    .dout19(r19tomtree0),
    .dout20(r20tomtree0),
    .dout21(r21tomtree0),
    .dout22(r22tomtree0),
    .dout23(r23tomtree0),
    .dout24(r24tomtree0),
    .dout25(r25tomtree0),
    .dout26(r26tomtree0),
    .dout27(r27tomtree0),
    .dout28(r28tomtree0),
    .dout29(r29tomtree0),
    .dout30(r30tomtree0),
    .dout31(r31tomtree0),
    .dout32(r32tomtree0),
    .dout33(r33tomtree0),
    .dout34(r34tomtree0),
    .dout35(r35tomtree0),
    .dout36(r36tomtree0),
    .dout37(r37tomtree0),
    .dout38(r38tomtree0),
    .dout39(r39tomtree0),
    .dout40(r40tomtree0),
    .dout41(r41tomtree0),
    .dout42(r42tomtree0),
    .dout43(r43tomtree0),
    .dout44(r44tomtree0),
    .dout45(r45tomtree0),
    .dout46(r46tomtree0),
    .dout47(r47tomtree0),
    .dout48(r48tomtree0),
    .dout49(r49tomtree0),
    .dout50(r50tomtree0),
    .dout51(r51tomtree0),
    .dout52(r52tomtree0),
    .dout53(r53tomtree0),
    .dout54(r54tomtree0),
    .dout55(r55tomtree0),
    .dout56(r56tomtree0),
    .dout57(r57tomtree0),
    .dout58(r58tomtree0),
    .dout59(r59tomtree0),
    .dout60(r60tomtree0),
    .dout61(r61tomtree0),
    .dout62(r62tomtree0),
    .dout63(r63tomtree0)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_1(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[1]),
    .din(mrgnsrcmuxout),
    .dout0(r64tomtree1),
    .dout1(r65tomtree1),
    .dout2(r66tomtree1),
    .dout3(r67tomtree1),
    .dout4(r68tomtree1),
    .dout5(r69tomtree1),
    .dout6(r70tomtree1),
    .dout7(r71tomtree1),
    .dout8(r72tomtree1),
    .dout9(r73tomtree1),
    .dout10(r74tomtree1),
    .dout11(r75tomtree1),
    .dout12(r76tomtree1),
    .dout13(r77tomtree1),
    .dout14(r78tomtree1),
    .dout15(r79tomtree1),
    .dout16(r80tomtree1),
    .dout17(r81tomtree1),
    .dout18(r82tomtree1),
    .dout19(r83tomtree1),
    .dout20(r84tomtree1),
    .dout21(r85tomtree1),
    .dout22(r86tomtree1),
    .dout23(r87tomtree1),
    .dout24(r88tomtree1),
    .dout25(r89tomtree1),
    .dout26(r90tomtree1),
    .dout27(r91tomtree1),
    .dout28(r92tomtree1),
    .dout29(r93tomtree1),
    .dout30(r94tomtree1),
    .dout31(r95tomtree1),
    .dout32(r96tomtree1),
    .dout33(r97tomtree1),
    .dout34(r98tomtree1),
    .dout35(r99tomtree1),
    .dout36(r100tomtree1),
    .dout37(r101tomtree1),
    .dout38(r102tomtree1),
    .dout39(r103tomtree1),
    .dout40(r104tomtree1),
    .dout41(r105tomtree1),
    .dout42(r106tomtree1),
    .dout43(r107tomtree1),
    .dout44(r108tomtree1),
    .dout45(r109tomtree1),
    .dout46(r110tomtree1),
    .dout47(r111tomtree1),
    .dout48(r112tomtree1),
    .dout49(r113tomtree1),
    .dout50(r114tomtree1),
    .dout51(r115tomtree1),
    .dout52(r116tomtree1),
    .dout53(r117tomtree1),
    .dout54(r118tomtree1),
    .dout55(r119tomtree1),
    .dout56(r120tomtree1),
    .dout57(r121tomtree1),
    .dout58(r122tomtree1),
    .dout59(r123tomtree1),
    .dout60(r124tomtree1),
    .dout61(r125tomtree1),
    .dout62(r126tomtree1),
    .dout63(r127tomtree1)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_2(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[2]),
    .din(mrgnsrcmuxout),
    .dout0(r128tomtree2),
    .dout1(r129tomtree2),
    .dout2(r130tomtree2),
    .dout3(r131tomtree2),
    .dout4(r132tomtree2),
    .dout5(r133tomtree2),
    .dout6(r134tomtree2),
    .dout7(r135tomtree2),
    .dout8(r136tomtree2),
    .dout9(r137tomtree2),
    .dout10(r138tomtree2),
    .dout11(r139tomtree2),
    .dout12(r140tomtree2),
    .dout13(r141tomtree2),
    .dout14(r142tomtree2),
    .dout15(r143tomtree2),
    .dout16(r144tomtree2),
    .dout17(r145tomtree2),
    .dout18(r146tomtree2),
    .dout19(r147tomtree2),
    .dout20(r148tomtree2),
    .dout21(r149tomtree2),
    .dout22(r150tomtree2),
    .dout23(r151tomtree2),
    .dout24(r152tomtree2),
    .dout25(r153tomtree2),
    .dout26(r154tomtree2),
    .dout27(r155tomtree2),
    .dout28(r156tomtree2),
    .dout29(r157tomtree2),
    .dout30(r158tomtree2),
    .dout31(r159tomtree2),
    .dout32(r160tomtree2),
    .dout33(r161tomtree2),
    .dout34(r162tomtree2),
    .dout35(r163tomtree2),
    .dout36(r164tomtree2),
    .dout37(r165tomtree2),
    .dout38(r166tomtree2),
    .dout39(r167tomtree2),
    .dout40(r168tomtree2),
    .dout41(r169tomtree2),
    .dout42(r170tomtree2),
    .dout43(r171tomtree2),
    .dout44(r172tomtree2),
    .dout45(r173tomtree2),
    .dout46(r174tomtree2),
    .dout47(r175tomtree2),
    .dout48(r176tomtree2),
    .dout49(r177tomtree2),
    .dout50(r178tomtree2),
    .dout51(r179tomtree2),
    .dout52(r180tomtree2),
    .dout53(r181tomtree2),
    .dout54(r182tomtree2),
    .dout55(r183tomtree2),
    .dout56(r184tomtree2),
    .dout57(r185tomtree2),
    .dout58(r186tomtree2),
    .dout59(r187tomtree2),
    .dout60(r188tomtree2),
    .dout61(r189tomtree2),
    .dout62(r190tomtree2),
    .dout63(r191tomtree2)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_3(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[3]),
    .din(mrgnsrcmuxout),
    .dout0(r192tomtree3),
    .dout1(r193tomtree3),
    .dout2(r194tomtree3),
    .dout3(r195tomtree3),
    .dout4(r196tomtree3),
    .dout5(r197tomtree3),
    .dout6(r198tomtree3),
    .dout7(r199tomtree3),
    .dout8(r200tomtree3),
    .dout9(r201tomtree3),
    .dout10(r202tomtree3),
    .dout11(r203tomtree3),
    .dout12(r204tomtree3),
    .dout13(r205tomtree3),
    .dout14(r206tomtree3),
    .dout15(r207tomtree3),
    .dout16(r208tomtree3),
    .dout17(r209tomtree3),
    .dout18(r210tomtree3),
    .dout19(r211tomtree3),
    .dout20(r212tomtree3),
    .dout21(r213tomtree3),
    .dout22(r214tomtree3),
    .dout23(r215tomtree3),
    .dout24(r216tomtree3),
    .dout25(r217tomtree3),
    .dout26(r218tomtree3),
    .dout27(r219tomtree3),
    .dout28(r220tomtree3),
    .dout29(r221tomtree3),
    .dout30(r222tomtree3),
    .dout31(r223tomtree3),
    .dout32(r224tomtree3),
    .dout33(r225tomtree3),
    .dout34(r226tomtree3),
    .dout35(r227tomtree3),
    .dout36(r228tomtree3),
    .dout37(r229tomtree3),
    .dout38(r230tomtree3),
    .dout39(r231tomtree3),
    .dout40(r232tomtree3),
    .dout41(r233tomtree3),
    .dout42(r234tomtree3),
    .dout43(r235tomtree3),
    .dout44(r236tomtree3),
    .dout45(r237tomtree3),
    .dout46(r238tomtree3),
    .dout47(r239tomtree3),
    .dout48(r240tomtree3),
    .dout49(r241tomtree3),
    .dout50(r242tomtree3),
    .dout51(r243tomtree3),
    .dout52(r244tomtree3),
    .dout53(r245tomtree3),
    .dout54(r246tomtree3),
    .dout55(r247tomtree3),
    .dout56(r248tomtree3),
    .dout57(r249tomtree3),
    .dout58(r250tomtree3),
    .dout59(r251tomtree3),
    .dout60(r252tomtree3),
    .dout61(r253tomtree3),
    .dout62(r254tomtree3),
    .dout63(r255tomtree3)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_4(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[4]),
    .din(mrgnsrcmuxout),
    .dout0(r256tomtree4),
    .dout1(r257tomtree4),
    .dout2(r258tomtree4),
    .dout3(r259tomtree4),
    .dout4(r260tomtree4),
    .dout5(r261tomtree4),
    .dout6(r262tomtree4),
    .dout7(r263tomtree4),
    .dout8(r264tomtree4),
    .dout9(r265tomtree4),
    .dout10(r266tomtree4),
    .dout11(r267tomtree4),
    .dout12(r268tomtree4),
    .dout13(r269tomtree4),
    .dout14(r270tomtree4),
    .dout15(r271tomtree4),
    .dout16(r272tomtree4),
    .dout17(r273tomtree4),
    .dout18(r274tomtree4),
    .dout19(r275tomtree4),
    .dout20(r276tomtree4),
    .dout21(r277tomtree4),
    .dout22(r278tomtree4),
    .dout23(r279tomtree4),
    .dout24(r280tomtree4),
    .dout25(r281tomtree4),
    .dout26(r282tomtree4),
    .dout27(r283tomtree4),
    .dout28(r284tomtree4),
    .dout29(r285tomtree4),
    .dout30(r286tomtree4),
    .dout31(r287tomtree4),
    .dout32(r288tomtree4),
    .dout33(r289tomtree4),
    .dout34(r290tomtree4),
    .dout35(r291tomtree4),
    .dout36(r292tomtree4),
    .dout37(r293tomtree4),
    .dout38(r294tomtree4),
    .dout39(r295tomtree4),
    .dout40(r296tomtree4),
    .dout41(r297tomtree4),
    .dout42(r298tomtree4),
    .dout43(r299tomtree4),
    .dout44(r300tomtree4),
    .dout45(r301tomtree4),
    .dout46(r302tomtree4),
    .dout47(r303tomtree4),
    .dout48(r304tomtree4),
    .dout49(r305tomtree4),
    .dout50(r306tomtree4),
    .dout51(r307tomtree4),
    .dout52(r308tomtree4),
    .dout53(r309tomtree4),
    .dout54(r310tomtree4),
    .dout55(r311tomtree4),
    .dout56(r312tomtree4),
    .dout57(r313tomtree4),
    .dout58(r314tomtree4),
    .dout59(r315tomtree4),
    .dout60(r316tomtree4),
    .dout61(r317tomtree4),
    .dout62(r318tomtree4),
    .dout63(r319tomtree4)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_5(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[5]),
    .din(mrgnsrcmuxout),
    .dout0(r320tomtree5),
    .dout1(r321tomtree5),
    .dout2(r322tomtree5),
    .dout3(r323tomtree5),
    .dout4(r324tomtree5),
    .dout5(r325tomtree5),
    .dout6(r326tomtree5),
    .dout7(r327tomtree5),
    .dout8(r328tomtree5),
    .dout9(r329tomtree5),
    .dout10(r330tomtree5),
    .dout11(r331tomtree5),
    .dout12(r332tomtree5),
    .dout13(r333tomtree5),
    .dout14(r334tomtree5),
    .dout15(r335tomtree5),
    .dout16(r336tomtree5),
    .dout17(r337tomtree5),
    .dout18(r338tomtree5),
    .dout19(r339tomtree5),
    .dout20(r340tomtree5),
    .dout21(r341tomtree5),
    .dout22(r342tomtree5),
    .dout23(r343tomtree5),
    .dout24(r344tomtree5),
    .dout25(r345tomtree5),
    .dout26(r346tomtree5),
    .dout27(r347tomtree5),
    .dout28(r348tomtree5),
    .dout29(r349tomtree5),
    .dout30(r350tomtree5),
    .dout31(r351tomtree5),
    .dout32(r352tomtree5),
    .dout33(r353tomtree5),
    .dout34(r354tomtree5),
    .dout35(r355tomtree5),
    .dout36(r356tomtree5),
    .dout37(r357tomtree5),
    .dout38(r358tomtree5),
    .dout39(r359tomtree5),
    .dout40(r360tomtree5),
    .dout41(r361tomtree5),
    .dout42(r362tomtree5),
    .dout43(r363tomtree5),
    .dout44(r364tomtree5),
    .dout45(r365tomtree5),
    .dout46(r366tomtree5),
    .dout47(r367tomtree5),
    .dout48(r368tomtree5),
    .dout49(r369tomtree5),
    .dout50(r370tomtree5),
    .dout51(r371tomtree5),
    .dout52(r372tomtree5),
    .dout53(r373tomtree5),
    .dout54(r374tomtree5),
    .dout55(r375tomtree5),
    .dout56(r376tomtree5),
    .dout57(r377tomtree5),
    .dout58(r378tomtree5),
    .dout59(r379tomtree5),
    .dout60(r380tomtree5),
    .dout61(r381tomtree5),
    .dout62(r382tomtree5),
    .dout63(r383tomtree5)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_6(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[6]),
    .din(mrgnsrcmuxout),
    .dout0(r384tomtree6),
    .dout1(r385tomtree6),
    .dout2(r386tomtree6),
    .dout3(r387tomtree6),
    .dout4(r388tomtree6),
    .dout5(r389tomtree6),
    .dout6(r390tomtree6),
    .dout7(r391tomtree6),
    .dout8(r392tomtree6),
    .dout9(r393tomtree6),
    .dout10(r394tomtree6),
    .dout11(r395tomtree6),
    .dout12(r396tomtree6),
    .dout13(r397tomtree6),
    .dout14(r398tomtree6),
    .dout15(r399tomtree6),
    .dout16(r400tomtree6),
    .dout17(r401tomtree6),
    .dout18(r402tomtree6),
    .dout19(r403tomtree6),
    .dout20(r404tomtree6),
    .dout21(r405tomtree6),
    .dout22(r406tomtree6),
    .dout23(r407tomtree6),
    .dout24(r408tomtree6),
    .dout25(r409tomtree6),
    .dout26(r410tomtree6),
    .dout27(r411tomtree6),
    .dout28(r412tomtree6),
    .dout29(r413tomtree6),
    .dout30(r414tomtree6),
    .dout31(r415tomtree6),
    .dout32(r416tomtree6),
    .dout33(r417tomtree6),
    .dout34(r418tomtree6),
    .dout35(r419tomtree6),
    .dout36(r420tomtree6),
    .dout37(r421tomtree6),
    .dout38(r422tomtree6),
    .dout39(r423tomtree6),
    .dout40(r424tomtree6),
    .dout41(r425tomtree6),
    .dout42(r426tomtree6),
    .dout43(r427tomtree6),
    .dout44(r428tomtree6),
    .dout45(r429tomtree6),
    .dout46(r430tomtree6),
    .dout47(r431tomtree6),
    .dout48(r432tomtree6),
    .dout49(r433tomtree6),
    .dout50(r434tomtree6),
    .dout51(r435tomtree6),
    .dout52(r436tomtree6),
    .dout53(r437tomtree6),
    .dout54(r438tomtree6),
    .dout55(r439tomtree6),
    .dout56(r440tomtree6),
    .dout57(r441tomtree6),
    .dout58(r442tomtree6),
    .dout59(r443tomtree6),
    .dout60(r444tomtree6),
    .dout61(r445tomtree6),
    .dout62(r446tomtree6),
    .dout63(r447tomtree6)
  );

  registers64 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RB_7(
    .clk(clk),
    .rst_n(rst_n),
    .en(rsrcmuxout),
    .cs(rbsrcmuxout[7]),
    .din(mrgnsrcmuxout),
    .dout0(r448tomtree7),
    .dout1(r449tomtree7),
    .dout2(r450tomtree7),
    .dout3(r451tomtree7),
    .dout4(r452tomtree7),
    .dout5(r453tomtree7),
    .dout6(r454tomtree7),
    .dout7(r455tomtree7),
    .dout8(r456tomtree7),
    .dout9(r457tomtree7),
    .dout10(r458tomtree7),
    .dout11(r459tomtree7),
    .dout12(r460tomtree7),
    .dout13(r461tomtree7),
    .dout14(r462tomtree7),
    .dout15(r463tomtree7),
    .dout16(r464tomtree7),
    .dout17(r465tomtree7),
    .dout18(r466tomtree7),
    .dout19(r467tomtree7),
    .dout20(r468tomtree7),
    .dout21(r469tomtree7),
    .dout22(r470tomtree7),
    .dout23(r471tomtree7),
    .dout24(r472tomtree7),
    .dout25(r473tomtree7),
    .dout26(r474tomtree7),
    .dout27(r475tomtree7),
    .dout28(r476tomtree7),
    .dout29(r477tomtree7),
    .dout30(r478tomtree7),
    .dout31(r479tomtree7),
    .dout32(r480tomtree7),
    .dout33(r481tomtree7),
    .dout34(r482tomtree7),
    .dout35(r483tomtree7),
    .dout36(r484tomtree7),
    .dout37(r485tomtree7),
    .dout38(r486tomtree7),
    .dout39(r487tomtree7),
    .dout40(r488tomtree7),
    .dout41(r489tomtree7),
    .dout42(r490tomtree7),
    .dout43(r491tomtree7),
    .dout44(r492tomtree7),
    .dout45(r493tomtree7),
    .dout46(r494tomtree7),
    .dout47(r495tomtree7),
    .dout48(r496tomtree7),
    .dout49(r497tomtree7),
    .dout50(r498tomtree7),
    .dout51(r499tomtree7),
    .dout52(r500tomtree7),
    .dout53(r501tomtree7),
    .dout54(r502tomtree7),
    .dout55(r503tomtree7),
    .dout56(r504tomtree7),
    .dout57(r505tomtree7),
    .dout58(r506tomtree7),
    .dout59(r507tomtree7),
    .dout60(r508tomtree7),
    .dout61(r509tomtree7),
    .dout62(r510tomtree7),
    .dout63(r511tomtree7)
  );
  
  mux2 #(.DATA_WIDTH(N_REGISTERSBANKS)) TrigMTreeSrcMux(
    .din0('b0), 
    .din1(decrb), 
    .sel(trigmtree), 
    .dout(trigmtreesrcmuxout)
  );
  
  register #(.DATA_WIDTH(N_REGISTERSBANKS)) RTrigMTreeSrcMux(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(trigmtreesrcmuxout),
    .dout(trigmtreeold)
  );
  
   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_0(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[0]),
    .din0(r0tomtree0),
    .din1(r1tomtree0),
    .din2(r2tomtree0),
    .din3(r3tomtree0),
    .din4(r4tomtree0),
    .din5(r5tomtree0),
    .din6(r6tomtree0),
    .din7(r7tomtree0),
    .din8(r8tomtree0),
    .din9(r9tomtree0),
    .din10(r10tomtree0),
    .din11(r11tomtree0),
    .din12(r12tomtree0),
    .din13(r13tomtree0),
    .din14(r14tomtree0),
    .din15(r15tomtree0),
    .din16(r16tomtree0),
    .din17(r17tomtree0),
    .din18(r18tomtree0),
    .din19(r19tomtree0),
    .din20(r20tomtree0),
    .din21(r21tomtree0),
    .din22(r22tomtree0),
    .din23(r23tomtree0),
    .din24(r24tomtree0),
    .din25(r25tomtree0),
    .din26(r26tomtree0),
    .din27(r27tomtree0),
    .din28(r28tomtree0),
    .din29(r29tomtree0),
    .din30(r30tomtree0),
    .din31(r31tomtree0),
    .din32(r32tomtree0),
    .din33(r33tomtree0),
    .din34(r34tomtree0),
    .din35(r35tomtree0),
    .din36(r36tomtree0),
    .din37(r37tomtree0),
    .din38(r38tomtree0),
    .din39(r39tomtree0),
    .din40(r40tomtree0),
    .din41(r41tomtree0),
    .din42(r42tomtree0),
    .din43(r43tomtree0),
    .din44(r44tomtree0),
    .din45(r45tomtree0),
    .din46(r46tomtree0),
    .din47(r47tomtree0),
    .din48(r48tomtree0),
    .din49(r49tomtree0),
    .din50(r50tomtree0),
    .din51(r51tomtree0),
    .din52(r52tomtree0),
    .din53(r53tomtree0),
    .din54(r54tomtree0),
    .din55(r55tomtree0),
    .din56(r56tomtree0),
    .din57(r57tomtree0),
    .din58(r58tomtree0),
    .din59(r59tomtree0),
    .din60(r60tomtree0),
    .din61(r61tomtree0),
    .din62(r62tomtree0),
    .din63(r63tomtree0),
    .max(mtree0tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_1(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[1]),
    .din0(r64tomtree1),
    .din1(r65tomtree1),
    .din2(r66tomtree1),
    .din3(r67tomtree1),
    .din4(r68tomtree1),
    .din5(r69tomtree1),
    .din6(r70tomtree1),
    .din7(r71tomtree1),
    .din8(r72tomtree1),
    .din9(r73tomtree1),
    .din10(r74tomtree1),
    .din11(r75tomtree1),
    .din12(r76tomtree1),
    .din13(r77tomtree1),
    .din14(r78tomtree1),
    .din15(r79tomtree1),
    .din16(r80tomtree1),
    .din17(r81tomtree1),
    .din18(r82tomtree1),
    .din19(r83tomtree1),
    .din20(r84tomtree1),
    .din21(r85tomtree1),
    .din22(r86tomtree1),
    .din23(r87tomtree1),
    .din24(r88tomtree1),
    .din25(r89tomtree1),
    .din26(r90tomtree1),
    .din27(r91tomtree1),
    .din28(r92tomtree1),
    .din29(r93tomtree1),
    .din30(r94tomtree1),
    .din31(r95tomtree1),
    .din32(r96tomtree1),
    .din33(r97tomtree1),
    .din34(r98tomtree1),
    .din35(r99tomtree1),
    .din36(r100tomtree1),
    .din37(r101tomtree1),
    .din38(r102tomtree1),
    .din39(r103tomtree1),
    .din40(r104tomtree1),
    .din41(r105tomtree1),
    .din42(r106tomtree1),
    .din43(r107tomtree1),
    .din44(r108tomtree1),
    .din45(r109tomtree1),
    .din46(r110tomtree1),
    .din47(r111tomtree1),
    .din48(r112tomtree1),
    .din49(r113tomtree1),
    .din50(r114tomtree1),
    .din51(r115tomtree1),
    .din52(r116tomtree1),
    .din53(r117tomtree1),
    .din54(r118tomtree1),
    .din55(r119tomtree1),
    .din56(r120tomtree1),
    .din57(r121tomtree1),
    .din58(r122tomtree1),
    .din59(r123tomtree1),
    .din60(r124tomtree1),
    .din61(r125tomtree1),
    .din62(r126tomtree1),
    .din63(r127tomtree1),
    .max(mtree1tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_2(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[2]),
    .din0(r128tomtree2),
    .din1(r129tomtree2),
    .din2(r130tomtree2),
    .din3(r131tomtree2),
    .din4(r132tomtree2),
    .din5(r133tomtree2),
    .din6(r134tomtree2),
    .din7(r135tomtree2),
    .din8(r136tomtree2),
    .din9(r137tomtree2),
    .din10(r138tomtree2),
    .din11(r139tomtree2),
    .din12(r140tomtree2),
    .din13(r141tomtree2),
    .din14(r142tomtree2),
    .din15(r143tomtree2),
    .din16(r144tomtree2),
    .din17(r145tomtree2),
    .din18(r146tomtree2),
    .din19(r147tomtree2),
    .din20(r148tomtree2),
    .din21(r149tomtree2),
    .din22(r150tomtree2),
    .din23(r151tomtree2),
    .din24(r152tomtree2),
    .din25(r153tomtree2),
    .din26(r154tomtree2),
    .din27(r155tomtree2),
    .din28(r156tomtree2),
    .din29(r157tomtree2),
    .din30(r158tomtree2),
    .din31(r159tomtree2),
    .din32(r160tomtree2),
    .din33(r161tomtree2),
    .din34(r162tomtree2),
    .din35(r163tomtree2),
    .din36(r164tomtree2),
    .din37(r165tomtree2),
    .din38(r166tomtree2),
    .din39(r167tomtree2),
    .din40(r168tomtree2),
    .din41(r169tomtree2),
    .din42(r170tomtree2),
    .din43(r171tomtree2),
    .din44(r172tomtree2),
    .din45(r173tomtree2),
    .din46(r174tomtree2),
    .din47(r175tomtree2),
    .din48(r176tomtree2),
    .din49(r177tomtree2),
    .din50(r178tomtree2),
    .din51(r179tomtree2),
    .din52(r180tomtree2),
    .din53(r181tomtree2),
    .din54(r182tomtree2),
    .din55(r183tomtree2),
    .din56(r184tomtree2),
    .din57(r185tomtree2),
    .din58(r186tomtree2),
    .din59(r187tomtree2),
    .din60(r188tomtree2),
    .din61(r189tomtree2),
    .din62(r190tomtree2),
    .din63(r191tomtree2),
    .max(mtree2tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_3(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[3]),
    .din0(r192tomtree3),
    .din1(r193tomtree3),
    .din2(r194tomtree3),
    .din3(r195tomtree3),
    .din4(r196tomtree3),
    .din5(r197tomtree3),
    .din6(r198tomtree3),
    .din7(r199tomtree3),
    .din8(r200tomtree3),
    .din9(r201tomtree3),
    .din10(r202tomtree3),
    .din11(r203tomtree3),
    .din12(r204tomtree3),
    .din13(r205tomtree3),
    .din14(r206tomtree3),
    .din15(r207tomtree3),
    .din16(r208tomtree3),
    .din17(r209tomtree3),
    .din18(r210tomtree3),
    .din19(r211tomtree3),
    .din20(r212tomtree3),
    .din21(r213tomtree3),
    .din22(r214tomtree3),
    .din23(r215tomtree3),
    .din24(r216tomtree3),
    .din25(r217tomtree3),
    .din26(r218tomtree3),
    .din27(r219tomtree3),
    .din28(r220tomtree3),
    .din29(r221tomtree3),
    .din30(r222tomtree3),
    .din31(r223tomtree3),
    .din32(r224tomtree3),
    .din33(r225tomtree3),
    .din34(r226tomtree3),
    .din35(r227tomtree3),
    .din36(r228tomtree3),
    .din37(r229tomtree3),
    .din38(r230tomtree3),
    .din39(r231tomtree3),
    .din40(r232tomtree3),
    .din41(r233tomtree3),
    .din42(r234tomtree3),
    .din43(r235tomtree3),
    .din44(r236tomtree3),
    .din45(r237tomtree3),
    .din46(r238tomtree3),
    .din47(r239tomtree3),
    .din48(r240tomtree3),
    .din49(r241tomtree3),
    .din50(r242tomtree3),
    .din51(r243tomtree3),
    .din52(r244tomtree3),
    .din53(r245tomtree3),
    .din54(r246tomtree3),
    .din55(r247tomtree3),
    .din56(r248tomtree3),
    .din57(r249tomtree3),
    .din58(r250tomtree3),
    .din59(r251tomtree3),
    .din60(r252tomtree3),
    .din61(r253tomtree3),
    .din62(r254tomtree3),
    .din63(r255tomtree3),
    .max(mtree3tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_4(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[4]),
    .din0(r256tomtree4),
    .din1(r257tomtree4),
    .din2(r258tomtree4),
    .din3(r259tomtree4),
    .din4(r260tomtree4),
    .din5(r261tomtree4),
    .din6(r262tomtree4),
    .din7(r263tomtree4),
    .din8(r264tomtree4),
    .din9(r265tomtree4),
    .din10(r266tomtree4),
    .din11(r267tomtree4),
    .din12(r268tomtree4),
    .din13(r269tomtree4),
    .din14(r270tomtree4),
    .din15(r271tomtree4),
    .din16(r272tomtree4),
    .din17(r273tomtree4),
    .din18(r274tomtree4),
    .din19(r275tomtree4),
    .din20(r276tomtree4),
    .din21(r277tomtree4),
    .din22(r278tomtree4),
    .din23(r279tomtree4),
    .din24(r280tomtree4),
    .din25(r281tomtree4),
    .din26(r282tomtree4),
    .din27(r283tomtree4),
    .din28(r284tomtree4),
    .din29(r285tomtree4),
    .din30(r286tomtree4),
    .din31(r287tomtree4),
    .din32(r288tomtree4),
    .din33(r289tomtree4),
    .din34(r290tomtree4),
    .din35(r291tomtree4),
    .din36(r292tomtree4),
    .din37(r293tomtree4),
    .din38(r294tomtree4),
    .din39(r295tomtree4),
    .din40(r296tomtree4),
    .din41(r297tomtree4),
    .din42(r298tomtree4),
    .din43(r299tomtree4),
    .din44(r300tomtree4),
    .din45(r301tomtree4),
    .din46(r302tomtree4),
    .din47(r303tomtree4),
    .din48(r304tomtree4),
    .din49(r305tomtree4),
    .din50(r306tomtree4),
    .din51(r307tomtree4),
    .din52(r308tomtree4),
    .din53(r309tomtree4),
    .din54(r310tomtree4),
    .din55(r311tomtree4),
    .din56(r312tomtree4),
    .din57(r313tomtree4),
    .din58(r314tomtree4),
    .din59(r315tomtree4),
    .din60(r316tomtree4),
    .din61(r317tomtree4),
    .din62(r318tomtree4),
    .din63(r319tomtree4),
    .max(mtree4tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_5(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[5]),
    .din0(r320tomtree5),
    .din1(r321tomtree5),
    .din2(r322tomtree5),
    .din3(r323tomtree5),
    .din4(r324tomtree5),
    .din5(r325tomtree5),
    .din6(r326tomtree5),
    .din7(r327tomtree5),
    .din8(r328tomtree5),
    .din9(r329tomtree5),
    .din10(r330tomtree5),
    .din11(r331tomtree5),
    .din12(r332tomtree5),
    .din13(r333tomtree5),
    .din14(r334tomtree5),
    .din15(r335tomtree5),
    .din16(r336tomtree5),
    .din17(r337tomtree5),
    .din18(r338tomtree5),
    .din19(r339tomtree5),
    .din20(r340tomtree5),
    .din21(r341tomtree5),
    .din22(r342tomtree5),
    .din23(r343tomtree5),
    .din24(r344tomtree5),
    .din25(r345tomtree5),
    .din26(r346tomtree5),
    .din27(r347tomtree5),
    .din28(r348tomtree5),
    .din29(r349tomtree5),
    .din30(r350tomtree5),
    .din31(r351tomtree5),
    .din32(r352tomtree5),
    .din33(r353tomtree5),
    .din34(r354tomtree5),
    .din35(r355tomtree5),
    .din36(r356tomtree5),
    .din37(r357tomtree5),
    .din38(r358tomtree5),
    .din39(r359tomtree5),
    .din40(r360tomtree5),
    .din41(r361tomtree5),
    .din42(r362tomtree5),
    .din43(r363tomtree5),
    .din44(r364tomtree5),
    .din45(r365tomtree5),
    .din46(r366tomtree5),
    .din47(r367tomtree5),
    .din48(r368tomtree5),
    .din49(r369tomtree5),
    .din50(r370tomtree5),
    .din51(r371tomtree5),
    .din52(r372tomtree5),
    .din53(r373tomtree5),
    .din54(r374tomtree5),
    .din55(r375tomtree5),
    .din56(r376tomtree5),
    .din57(r377tomtree5),
    .din58(r378tomtree5),
    .din59(r379tomtree5),
    .din60(r380tomtree5),
    .din61(r381tomtree5),
    .din62(r382tomtree5),
    .din63(r383tomtree5),
    .max(mtree5tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_6(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[6]),
    .din0(r384tomtree6),
    .din1(r385tomtree6),
    .din2(r386tomtree6),
    .din3(r387tomtree6),
    .din4(r388tomtree6),
    .din5(r389tomtree6),
    .din6(r390tomtree6),
    .din7(r391tomtree6),
    .din8(r392tomtree6),
    .din9(r393tomtree6),
    .din10(r394tomtree6),
    .din11(r395tomtree6),
    .din12(r396tomtree6),
    .din13(r397tomtree6),
    .din14(r398tomtree6),
    .din15(r399tomtree6),
    .din16(r400tomtree6),
    .din17(r401tomtree6),
    .din18(r402tomtree6),
    .din19(r403tomtree6),
    .din20(r404tomtree6),
    .din21(r405tomtree6),
    .din22(r406tomtree6),
    .din23(r407tomtree6),
    .din24(r408tomtree6),
    .din25(r409tomtree6),
    .din26(r410tomtree6),
    .din27(r411tomtree6),
    .din28(r412tomtree6),
    .din29(r413tomtree6),
    .din30(r414tomtree6),
    .din31(r415tomtree6),
    .din32(r416tomtree6),
    .din33(r417tomtree6),
    .din34(r418tomtree6),
    .din35(r419tomtree6),
    .din36(r420tomtree6),
    .din37(r421tomtree6),
    .din38(r422tomtree6),
    .din39(r423tomtree6),
    .din40(r424tomtree6),
    .din41(r425tomtree6),
    .din42(r426tomtree6),
    .din43(r427tomtree6),
    .din44(r428tomtree6),
    .din45(r429tomtree6),
    .din46(r430tomtree6),
    .din47(r431tomtree6),
    .din48(r432tomtree6),
    .din49(r433tomtree6),
    .din50(r434tomtree6),
    .din51(r435tomtree6),
    .din52(r436tomtree6),
    .din53(r437tomtree6),
    .din54(r438tomtree6),
    .din55(r439tomtree6),
    .din56(r440tomtree6),
    .din57(r441tomtree6),
    .din58(r442tomtree6),
    .din59(r443tomtree6),
    .din60(r444tomtree6),
    .din61(r445tomtree6),
    .din62(r446tomtree6),
    .din63(r447tomtree6),
    .max(mtree6tomaxsrcmux)
  );

   maxtree64 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) MTree_7(
    .clk(clk),
    .rst_n(rst_n),
    .start(1'b1),//.start(trigmtreeold[7]),
    .din0(r448tomtree7),
    .din1(r449tomtree7),
    .din2(r450tomtree7),
    .din3(r451tomtree7),
    .din4(r452tomtree7),
    .din5(r453tomtree7),
    .din6(r454tomtree7),
    .din7(r455tomtree7),
    .din8(r456tomtree7),
    .din9(r457tomtree7),
    .din10(r458tomtree7),
    .din11(r459tomtree7),
    .din12(r460tomtree7),
    .din13(r461tomtree7),
    .din14(r462tomtree7),
    .din15(r463tomtree7),
    .din16(r464tomtree7),
    .din17(r465tomtree7),
    .din18(r466tomtree7),
    .din19(r467tomtree7),
    .din20(r468tomtree7),
    .din21(r469tomtree7),
    .din22(r470tomtree7),
    .din23(r471tomtree7),
    .din24(r472tomtree7),
    .din25(r473tomtree7),
    .din26(r474tomtree7),
    .din27(r475tomtree7),
    .din28(r476tomtree7),
    .din29(r477tomtree7),
    .din30(r478tomtree7),
    .din31(r479tomtree7),
    .din32(r480tomtree7),
    .din33(r481tomtree7),
    .din34(r482tomtree7),
    .din35(r483tomtree7),
    .din36(r484tomtree7),
    .din37(r485tomtree7),
    .din38(r486tomtree7),
    .din39(r487tomtree7),
    .din40(r488tomtree7),
    .din41(r489tomtree7),
    .din42(r490tomtree7),
    .din43(r491tomtree7),
    .din44(r492tomtree7),
    .din45(r493tomtree7),
    .din46(r494tomtree7),
    .din47(r495tomtree7),
    .din48(r496tomtree7),
    .din49(r497tomtree7),
    .din50(r498tomtree7),
    .din51(r499tomtree7),
    .din52(r500tomtree7),
    .din53(r501tomtree7),
    .din54(r502tomtree7),
    .din55(r503tomtree7),
    .din56(r504tomtree7),
    .din57(r505tomtree7),
    .din58(r506tomtree7),
    .din59(r507tomtree7),
    .din60(r508tomtree7),
    .din61(r509tomtree7),
    .din62(r510tomtree7),
    .din63(r511tomtree7),
    .max(mtree7tomaxsrcmux)
  );
  
  mux8 #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) MaxSrcMux(
    .din0(mtree0tomaxsrcmux),
    .din1(mtree1tomaxsrcmux),
    .din2(mtree2tomaxsrcmux),
    .din3(mtree3tomaxsrcmux),
    .din4(mtree4tomaxsrcmux),
    .din5(mtree5tomaxsrcmux),
    .din6(mtree6tomaxsrcmux),
    .din7(mtree7tomaxsrcmux),
    .sel(rcntrb),
    .dout(maxsrcmuxtocmp)
  );

  comparator #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH), .N_REGISTERS(N_REGISTERS)) Cmp(
    .max(maxsrcmuxtocmp),
    .margin({mrgnindx,mrgn}),
    .trig(trigmax),
    .r_sel(rcmp),
    .dout(mrgncmp)
  );
  
  register #(.DATA_WIDTH(1)) RCmpTrig(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(trigmax),
    .dout(rtrigmax)
  );
  
  register #(.DATA_WIDTH($clog2(N_REGISTERS))) RCmpRSel(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(rcmp),
    .dout(rrcmp)
  );
  
  register #(.DATA_WIDTH(DATA_WIDTH+INDX_WIDTH+ADDR_WIDTH)) RCmpMrgn(
    .clk(clk),
    .rst_n(rst_n),
    .en(1'b1),
    .cs(1'b1),
    .din(mrgncmp),
    .dout(rmrgncmp)
  );
  
  mux512 #(.DATA_WIDTH(DATA_WIDTH), .INDX_WIDTH(INDX_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) OutSrcMux(
    .din0(r0tomtree0),
    .din1(r1tomtree0),
    .din2(r2tomtree0),
    .din3(r3tomtree0),
    .din4(r4tomtree0),
    .din5(r5tomtree0),
    .din6(r6tomtree0),
    .din7(r7tomtree0),
    .din8(r8tomtree0),
    .din9(r9tomtree0),
    .din10(r10tomtree0),
    .din11(r11tomtree0),
    .din12(r12tomtree0),
    .din13(r13tomtree0),
    .din14(r14tomtree0),
    .din15(r15tomtree0),
    .din16(r16tomtree0),
    .din17(r17tomtree0),
    .din18(r18tomtree0),
    .din19(r19tomtree0),
    .din20(r20tomtree0),
    .din21(r21tomtree0),
    .din22(r22tomtree0),
    .din23(r23tomtree0),
    .din24(r24tomtree0),
    .din25(r25tomtree0),
    .din26(r26tomtree0),
    .din27(r27tomtree0),
    .din28(r28tomtree0),
    .din29(r29tomtree0),
    .din30(r30tomtree0),
    .din31(r31tomtree0),
    .din32(r32tomtree0),
    .din33(r33tomtree0),
    .din34(r34tomtree0),
    .din35(r35tomtree0),
    .din36(r36tomtree0),
    .din37(r37tomtree0),
    .din38(r38tomtree0),
    .din39(r39tomtree0),
    .din40(r40tomtree0),
    .din41(r41tomtree0),
    .din42(r42tomtree0),
    .din43(r43tomtree0),
    .din44(r44tomtree0),
    .din45(r45tomtree0),
    .din46(r46tomtree0),
    .din47(r47tomtree0),
    .din48(r48tomtree0),
    .din49(r49tomtree0),
    .din50(r50tomtree0),
    .din51(r51tomtree0),
    .din52(r52tomtree0),
    .din53(r53tomtree0),
    .din54(r54tomtree0),
    .din55(r55tomtree0),
    .din56(r56tomtree0),
    .din57(r57tomtree0),
    .din58(r58tomtree0),
    .din59(r59tomtree0),
    .din60(r60tomtree0),
    .din61(r61tomtree0),
    .din62(r62tomtree0),
    .din63(r63tomtree0),
    .din64(r64tomtree1),
    .din65(r65tomtree1),
    .din66(r66tomtree1),
    .din67(r67tomtree1),
    .din68(r68tomtree1),
    .din69(r69tomtree1),
    .din70(r70tomtree1),
    .din71(r71tomtree1),
    .din72(r72tomtree1),
    .din73(r73tomtree1),
    .din74(r74tomtree1),
    .din75(r75tomtree1),
    .din76(r76tomtree1),
    .din77(r77tomtree1),
    .din78(r78tomtree1),
    .din79(r79tomtree1),
    .din80(r80tomtree1),
    .din81(r81tomtree1),
    .din82(r82tomtree1),
    .din83(r83tomtree1),
    .din84(r84tomtree1),
    .din85(r85tomtree1),
    .din86(r86tomtree1),
    .din87(r87tomtree1),
    .din88(r88tomtree1),
    .din89(r89tomtree1),
    .din90(r90tomtree1),
    .din91(r91tomtree1),
    .din92(r92tomtree1),
    .din93(r93tomtree1),
    .din94(r94tomtree1),
    .din95(r95tomtree1),
    .din96(r96tomtree1),
    .din97(r97tomtree1),
    .din98(r98tomtree1),
    .din99(r99tomtree1),
    .din100(r100tomtree1),
    .din101(r101tomtree1),
    .din102(r102tomtree1),
    .din103(r103tomtree1),
    .din104(r104tomtree1),
    .din105(r105tomtree1),
    .din106(r106tomtree1),
    .din107(r107tomtree1),
    .din108(r108tomtree1),
    .din109(r109tomtree1),
    .din110(r110tomtree1),
    .din111(r111tomtree1),
    .din112(r112tomtree1),
    .din113(r113tomtree1),
    .din114(r114tomtree1),
    .din115(r115tomtree1),
    .din116(r116tomtree1),
    .din117(r117tomtree1),
    .din118(r118tomtree1),
    .din119(r119tomtree1),
    .din120(r120tomtree1),
    .din121(r121tomtree1),
    .din122(r122tomtree1),
    .din123(r123tomtree1),
    .din124(r124tomtree1),
    .din125(r125tomtree1),
    .din126(r126tomtree1),
    .din127(r127tomtree1),
    .din128(r128tomtree2),
    .din129(r129tomtree2),
    .din130(r130tomtree2),
    .din131(r131tomtree2),
    .din132(r132tomtree2),
    .din133(r133tomtree2),
    .din134(r134tomtree2),
    .din135(r135tomtree2),
    .din136(r136tomtree2),
    .din137(r137tomtree2),
    .din138(r138tomtree2),
    .din139(r139tomtree2),
    .din140(r140tomtree2),
    .din141(r141tomtree2),
    .din142(r142tomtree2),
    .din143(r143tomtree2),
    .din144(r144tomtree2),
    .din145(r145tomtree2),
    .din146(r146tomtree2),
    .din147(r147tomtree2),
    .din148(r148tomtree2),
    .din149(r149tomtree2),
    .din150(r150tomtree2),
    .din151(r151tomtree2),
    .din152(r152tomtree2),
    .din153(r153tomtree2),
    .din154(r154tomtree2),
    .din155(r155tomtree2),
    .din156(r156tomtree2),
    .din157(r157tomtree2),
    .din158(r158tomtree2),
    .din159(r159tomtree2),
    .din160(r160tomtree2),
    .din161(r161tomtree2),
    .din162(r162tomtree2),
    .din163(r163tomtree2),
    .din164(r164tomtree2),
    .din165(r165tomtree2),
    .din166(r166tomtree2),
    .din167(r167tomtree2),
    .din168(r168tomtree2),
    .din169(r169tomtree2),
    .din170(r170tomtree2),
    .din171(r171tomtree2),
    .din172(r172tomtree2),
    .din173(r173tomtree2),
    .din174(r174tomtree2),
    .din175(r175tomtree2),
    .din176(r176tomtree2),
    .din177(r177tomtree2),
    .din178(r178tomtree2),
    .din179(r179tomtree2),
    .din180(r180tomtree2),
    .din181(r181tomtree2),
    .din182(r182tomtree2),
    .din183(r183tomtree2),
    .din184(r184tomtree2),
    .din185(r185tomtree2),
    .din186(r186tomtree2),
    .din187(r187tomtree2),
    .din188(r188tomtree2),
    .din189(r189tomtree2),
    .din190(r190tomtree2),
    .din191(r191tomtree2),
    .din192(r192tomtree3),
    .din193(r193tomtree3),
    .din194(r194tomtree3),
    .din195(r195tomtree3),
    .din196(r196tomtree3),
    .din197(r197tomtree3),
    .din198(r198tomtree3),
    .din199(r199tomtree3),
    .din200(r200tomtree3),
    .din201(r201tomtree3),
    .din202(r202tomtree3),
    .din203(r203tomtree3),
    .din204(r204tomtree3),
    .din205(r205tomtree3),
    .din206(r206tomtree3),
    .din207(r207tomtree3),
    .din208(r208tomtree3),
    .din209(r209tomtree3),
    .din210(r210tomtree3),
    .din211(r211tomtree3),
    .din212(r212tomtree3),
    .din213(r213tomtree3),
    .din214(r214tomtree3),
    .din215(r215tomtree3),
    .din216(r216tomtree3),
    .din217(r217tomtree3),
    .din218(r218tomtree3),
    .din219(r219tomtree3),
    .din220(r220tomtree3),
    .din221(r221tomtree3),
    .din222(r222tomtree3),
    .din223(r223tomtree3),
    .din224(r224tomtree3),
    .din225(r225tomtree3),
    .din226(r226tomtree3),
    .din227(r227tomtree3),
    .din228(r228tomtree3),
    .din229(r229tomtree3),
    .din230(r230tomtree3),
    .din231(r231tomtree3),
    .din232(r232tomtree3),
    .din233(r233tomtree3),
    .din234(r234tomtree3),
    .din235(r235tomtree3),
    .din236(r236tomtree3),
    .din237(r237tomtree3),
    .din238(r238tomtree3),
    .din239(r239tomtree3),
    .din240(r240tomtree3),
    .din241(r241tomtree3),
    .din242(r242tomtree3),
    .din243(r243tomtree3),
    .din244(r244tomtree3),
    .din245(r245tomtree3),
    .din246(r246tomtree3),
    .din247(r247tomtree3),
    .din248(r248tomtree3),
    .din249(r249tomtree3),
    .din250(r250tomtree3),
    .din251(r251tomtree3),
    .din252(r252tomtree3),
    .din253(r253tomtree3),
    .din254(r254tomtree3),
    .din255(r255tomtree3),
    .din256(r256tomtree4),
    .din257(r257tomtree4),
    .din258(r258tomtree4),
    .din259(r259tomtree4),
    .din260(r260tomtree4),
    .din261(r261tomtree4),
    .din262(r262tomtree4),
    .din263(r263tomtree4),
    .din264(r264tomtree4),
    .din265(r265tomtree4),
    .din266(r266tomtree4),
    .din267(r267tomtree4),
    .din268(r268tomtree4),
    .din269(r269tomtree4),
    .din270(r270tomtree4),
    .din271(r271tomtree4),
    .din272(r272tomtree4),
    .din273(r273tomtree4),
    .din274(r274tomtree4),
    .din275(r275tomtree4),
    .din276(r276tomtree4),
    .din277(r277tomtree4),
    .din278(r278tomtree4),
    .din279(r279tomtree4),
    .din280(r280tomtree4),
    .din281(r281tomtree4),
    .din282(r282tomtree4),
    .din283(r283tomtree4),
    .din284(r284tomtree4),
    .din285(r285tomtree4),
    .din286(r286tomtree4),
    .din287(r287tomtree4),
    .din288(r288tomtree4),
    .din289(r289tomtree4),
    .din290(r290tomtree4),
    .din291(r291tomtree4),
    .din292(r292tomtree4),
    .din293(r293tomtree4),
    .din294(r294tomtree4),
    .din295(r295tomtree4),
    .din296(r296tomtree4),
    .din297(r297tomtree4),
    .din298(r298tomtree4),
    .din299(r299tomtree4),
    .din300(r300tomtree4),
    .din301(r301tomtree4),
    .din302(r302tomtree4),
    .din303(r303tomtree4),
    .din304(r304tomtree4),
    .din305(r305tomtree4),
    .din306(r306tomtree4),
    .din307(r307tomtree4),
    .din308(r308tomtree4),
    .din309(r309tomtree4),
    .din310(r310tomtree4),
    .din311(r311tomtree4),
    .din312(r312tomtree4),
    .din313(r313tomtree4),
    .din314(r314tomtree4),
    .din315(r315tomtree4),
    .din316(r316tomtree4),
    .din317(r317tomtree4),
    .din318(r318tomtree4),
    .din319(r319tomtree4),
    .din320(r320tomtree5),
    .din321(r321tomtree5),
    .din322(r322tomtree5),
    .din323(r323tomtree5),
    .din324(r324tomtree5),
    .din325(r325tomtree5),
    .din326(r326tomtree5),
    .din327(r327tomtree5),
    .din328(r328tomtree5),
    .din329(r329tomtree5),
    .din330(r330tomtree5),
    .din331(r331tomtree5),
    .din332(r332tomtree5),
    .din333(r333tomtree5),
    .din334(r334tomtree5),
    .din335(r335tomtree5),
    .din336(r336tomtree5),
    .din337(r337tomtree5),
    .din338(r338tomtree5),
    .din339(r339tomtree5),
    .din340(r340tomtree5),
    .din341(r341tomtree5),
    .din342(r342tomtree5),
    .din343(r343tomtree5),
    .din344(r344tomtree5),
    .din345(r345tomtree5),
    .din346(r346tomtree5),
    .din347(r347tomtree5),
    .din348(r348tomtree5),
    .din349(r349tomtree5),
    .din350(r350tomtree5),
    .din351(r351tomtree5),
    .din352(r352tomtree5),
    .din353(r353tomtree5),
    .din354(r354tomtree5),
    .din355(r355tomtree5),
    .din356(r356tomtree5),
    .din357(r357tomtree5),
    .din358(r358tomtree5),
    .din359(r359tomtree5),
    .din360(r360tomtree5),
    .din361(r361tomtree5),
    .din362(r362tomtree5),
    .din363(r363tomtree5),
    .din364(r364tomtree5),
    .din365(r365tomtree5),
    .din366(r366tomtree5),
    .din367(r367tomtree5),
    .din368(r368tomtree5),
    .din369(r369tomtree5),
    .din370(r370tomtree5),
    .din371(r371tomtree5),
    .din372(r372tomtree5),
    .din373(r373tomtree5),
    .din374(r374tomtree5),
    .din375(r375tomtree5),
    .din376(r376tomtree5),
    .din377(r377tomtree5),
    .din378(r378tomtree5),
    .din379(r379tomtree5),
    .din380(r380tomtree5),
    .din381(r381tomtree5),
    .din382(r382tomtree5),
    .din383(r383tomtree5),
    .din384(r384tomtree6),
    .din385(r385tomtree6),
    .din386(r386tomtree6),
    .din387(r387tomtree6),
    .din388(r388tomtree6),
    .din389(r389tomtree6),
    .din390(r390tomtree6),
    .din391(r391tomtree6),
    .din392(r392tomtree6),
    .din393(r393tomtree6),
    .din394(r394tomtree6),
    .din395(r395tomtree6),
    .din396(r396tomtree6),
    .din397(r397tomtree6),
    .din398(r398tomtree6),
    .din399(r399tomtree6),
    .din400(r400tomtree6),
    .din401(r401tomtree6),
    .din402(r402tomtree6),
    .din403(r403tomtree6),
    .din404(r404tomtree6),
    .din405(r405tomtree6),
    .din406(r406tomtree6),
    .din407(r407tomtree6),
    .din408(r408tomtree6),
    .din409(r409tomtree6),
    .din410(r410tomtree6),
    .din411(r411tomtree6),
    .din412(r412tomtree6),
    .din413(r413tomtree6),
    .din414(r414tomtree6),
    .din415(r415tomtree6),
    .din416(r416tomtree6),
    .din417(r417tomtree6),
    .din418(r418tomtree6),
    .din419(r419tomtree6),
    .din420(r420tomtree6),
    .din421(r421tomtree6),
    .din422(r422tomtree6),
    .din423(r423tomtree6),
    .din424(r424tomtree6),
    .din425(r425tomtree6),
    .din426(r426tomtree6),
    .din427(r427tomtree6),
    .din428(r428tomtree6),
    .din429(r429tomtree6),
    .din430(r430tomtree6),
    .din431(r431tomtree6),
    .din432(r432tomtree6),
    .din433(r433tomtree6),
    .din434(r434tomtree6),
    .din435(r435tomtree6),
    .din436(r436tomtree6),
    .din437(r437tomtree6),
    .din438(r438tomtree6),
    .din439(r439tomtree6),
    .din440(r440tomtree6),
    .din441(r441tomtree6),
    .din442(r442tomtree6),
    .din443(r443tomtree6),
    .din444(r444tomtree6),
    .din445(r445tomtree6),
    .din446(r446tomtree6),
    .din447(r447tomtree6),
    .din448(r448tomtree7),
    .din449(r449tomtree7),
    .din450(r450tomtree7),
    .din451(r451tomtree7),
    .din452(r452tomtree7),
    .din453(r453tomtree7),
    .din454(r454tomtree7),
    .din455(r455tomtree7),
    .din456(r456tomtree7),
    .din457(r457tomtree7),
    .din458(r458tomtree7),
    .din459(r459tomtree7),
    .din460(r460tomtree7),
    .din461(r461tomtree7),
    .din462(r462tomtree7),
    .din463(r463tomtree7),
    .din464(r464tomtree7),
    .din465(r465tomtree7),
    .din466(r466tomtree7),
    .din467(r467tomtree7),
    .din468(r468tomtree7),
    .din469(r469tomtree7),
    .din470(r470tomtree7),
    .din471(r471tomtree7),
    .din472(r472tomtree7),
    .din473(r473tomtree7),
    .din474(r474tomtree7),
    .din475(r475tomtree7),
    .din476(r476tomtree7),
    .din477(r477tomtree7),
    .din478(r478tomtree7),
    .din479(r479tomtree7),
    .din480(r480tomtree7),
    .din481(r481tomtree7),
    .din482(r482tomtree7),
    .din483(r483tomtree7),
    .din484(r484tomtree7),
    .din485(r485tomtree7),
    .din486(r486tomtree7),
    .din487(r487tomtree7),
    .din488(r488tomtree7),
    .din489(r489tomtree7),
    .din490(r490tomtree7),
    .din491(r491tomtree7),
    .din492(r492tomtree7),
    .din493(r493tomtree7),
    .din494(r494tomtree7),
    .din495(r495tomtree7),
    .din496(r496tomtree7),
    .din497(r497tomtree7),
    .din498(r498tomtree7),
    .din499(r499tomtree7),
    .din500(r500tomtree7),
    .din501(r501tomtree7),
    .din502(r502tomtree7),
    .din503(r503tomtree7),
    .din504(r504tomtree7),
    .din505(r505tomtree7),
    .din506(r506tomtree7),
    .din507(r507tomtree7),
    .din508(r508tomtree7),
    .din509(r509tomtree7),
    .din510(r510tomtree7),
    .din511(r511tomtree7),
    .sel(cntout),
    .indx(indx)
  );

  counter_out #(.INCR(1), .CNT_WIDTH($clog2(BATCH_SIZE))) CntOut(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntouten),
    .cnt(cntout)
  );

  counter_addr #(.INCR(ADDR_INCR_PORTB), .ADDR_WIDTH(ADDR_WIDTH_PORTB)) CntAddrB(
    .clk(clk),
    .rst_n(rst_n),
    .en(cntaddrben),
    .cnt(addrbw)
  );
  
  //bram output port
  assign clkb = clk;
  assign rstb = ~rst_n;
  assign enb = enbw;
  assign addrb = addrbw;
  assign dinb = indx;
  assign web = webw;
  
endmodule